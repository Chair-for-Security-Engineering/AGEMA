
module SkinnyTop_GHPC_ANF_ClockGating_d1 ( Plaintext_s0, Key_s0, clk, rst, 
        Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch
 );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Plaintext_s1;
  input [63:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  input clk, rst;
  output done, Synch;
  wire   signal_1166, signal_1099, signal_1164, signal_1163, signal_1169,
         signal_1098, signal_1167, signal_1162, signal_1172, signal_1097,
         signal_1170, signal_1161, signal_1175, signal_1096, signal_1173,
         signal_1160, signal_1178, signal_1095, signal_1176, signal_1159,
         signal_1181, signal_1094, signal_1179, signal_1158, signal_1184,
         signal_1093, signal_1182, signal_1157, signal_1187, signal_1092,
         signal_1185, signal_1156, signal_1190, signal_1091, signal_1188,
         signal_1155, signal_1193, signal_1090, signal_1191, signal_1154,
         signal_1196, signal_1089, signal_1194, signal_1153, signal_1199,
         signal_1088, signal_1197, signal_1152, signal_1202, signal_1087,
         signal_1200, signal_1151, signal_1205, signal_1086, signal_1203,
         signal_1150, signal_1208, signal_1085, signal_1206, signal_1149,
         signal_1211, signal_1084, signal_1209, signal_1148, signal_1214,
         signal_1083, signal_1212, signal_1147, signal_1217, signal_1082,
         signal_1215, signal_1146, signal_1220, signal_1081, signal_1218,
         signal_1145, signal_1223, signal_1080, signal_1221, signal_1144,
         signal_1226, signal_1079, signal_1224, signal_1143, signal_1229,
         signal_1078, signal_1227, signal_1142, signal_1232, signal_1077,
         signal_1230, signal_1141, signal_1235, signal_1076, signal_1233,
         signal_1140, signal_1238, signal_1075, signal_1236, signal_1139,
         signal_1241, signal_1074, signal_1239, signal_1138, signal_1244,
         signal_1073, signal_1242, signal_1137, signal_1247, signal_1072,
         signal_1245, signal_1136, signal_1250, signal_1071, signal_1248,
         signal_1135, signal_1253, signal_1070, signal_1251, signal_1134,
         signal_1256, signal_1069, signal_1254, signal_1133, signal_1259,
         signal_1068, signal_1257, signal_1132, signal_1262, signal_1067,
         signal_1260, signal_1131, signal_1265, signal_1066, signal_1263,
         signal_1130, signal_1268, signal_1065, signal_1266, signal_1129,
         signal_1271, signal_1064, signal_1269, signal_1128, signal_1274,
         signal_1063, signal_1272, signal_1127, signal_1277, signal_1062,
         signal_1275, signal_1126, signal_1280, signal_1061, signal_1278,
         signal_1125, signal_1283, signal_1060, signal_1281, signal_1124,
         signal_1286, signal_1059, signal_1284, signal_1123, signal_1289,
         signal_1058, signal_1287, signal_1122, signal_1292, signal_1057,
         signal_1290, signal_1121, signal_1295, signal_1056, signal_1293,
         signal_1120, signal_1298, signal_1055, signal_1296, signal_1119,
         signal_1301, signal_1054, signal_1299, signal_1118, signal_1304,
         signal_1053, signal_1302, signal_1117, signal_1307, signal_1052,
         signal_1305, signal_1116, signal_1310, signal_1051, signal_1308,
         signal_1115, signal_1313, signal_1050, signal_1311, signal_1114,
         signal_1316, signal_1049, signal_1314, signal_1113, signal_1319,
         signal_1048, signal_1317, signal_1112, signal_1322, signal_1047,
         signal_1320, signal_1111, signal_1325, signal_1046, signal_1323,
         signal_1110, signal_1328, signal_1045, signal_1326, signal_1109,
         signal_1331, signal_1044, signal_1329, signal_1108, signal_1334,
         signal_1043, signal_1332, signal_1107, signal_1337, signal_1042,
         signal_1335, signal_1106, signal_1340, signal_1041, signal_1338,
         signal_1105, signal_1343, signal_1040, signal_1341, signal_1104,
         signal_1346, signal_1039, signal_1344, signal_1103, signal_1349,
         signal_1038, signal_1347, signal_1102, signal_1352, signal_1037,
         signal_1350, signal_1101, signal_1355, signal_1036, signal_1353,
         signal_1100, signal_1035, signal_1028, signal_1034, signal_1033,
         signal_1026, signal_1032, signal_1025, signal_1031, signal_1030,
         signal_940, signal_939, signal_943, signal_1676, signal_1485,
         signal_903, signal_1483, signal_839, signal_1487, signal_902,
         signal_1482, signal_838, signal_1489, signal_901, signal_1481,
         signal_837, signal_1491, signal_900, signal_1480, signal_836,
         signal_1493, signal_899, signal_1479, signal_835, signal_1495,
         signal_898, signal_1478, signal_834, signal_1497, signal_897,
         signal_1477, signal_833, signal_1499, signal_896, signal_1476,
         signal_832, signal_1501, signal_895, signal_1475, signal_831,
         signal_1503, signal_894, signal_1474, signal_830, signal_1505,
         signal_893, signal_1473, signal_829, signal_1507, signal_892,
         signal_1472, signal_828, signal_1509, signal_891, signal_1471,
         signal_827, signal_1511, signal_890, signal_1470, signal_826,
         signal_1513, signal_889, signal_1469, signal_825, signal_1515,
         signal_888, signal_1468, signal_824, signal_1517, signal_887,
         signal_1467, signal_823, signal_1519, signal_886, signal_1466,
         signal_822, signal_1521, signal_885, signal_1465, signal_821,
         signal_1523, signal_884, signal_1464, signal_820, signal_1525,
         signal_883, signal_1463, signal_819, signal_1527, signal_882,
         signal_1462, signal_818, signal_1529, signal_881, signal_1461,
         signal_817, signal_1531, signal_880, signal_1460, signal_816,
         signal_1533, signal_879, signal_1459, signal_815, signal_1535,
         signal_878, signal_1458, signal_814, signal_1537, signal_877,
         signal_1457, signal_813, signal_1539, signal_876, signal_1456,
         signal_812, signal_1541, signal_875, signal_1455, signal_811,
         signal_1543, signal_874, signal_1454, signal_810, signal_1545,
         signal_873, signal_1453, signal_809, signal_1547, signal_872,
         signal_1452, signal_808, signal_1549, signal_871, signal_1451,
         signal_807, signal_1551, signal_870, signal_1450, signal_806,
         signal_1553, signal_869, signal_1449, signal_805, signal_1555,
         signal_868, signal_1448, signal_804, signal_1557, signal_867,
         signal_1447, signal_803, signal_1559, signal_866, signal_1446,
         signal_802, signal_1561, signal_865, signal_1445, signal_801,
         signal_1563, signal_864, signal_1444, signal_800, signal_1565,
         signal_863, signal_1443, signal_799, signal_1567, signal_862,
         signal_1442, signal_798, signal_1569, signal_861, signal_1441,
         signal_797, signal_1571, signal_860, signal_1440, signal_796,
         signal_1573, signal_859, signal_1439, signal_795, signal_1575,
         signal_858, signal_1438, signal_794, signal_1577, signal_857,
         signal_1437, signal_793, signal_1579, signal_856, signal_1436,
         signal_792, signal_1581, signal_855, signal_1435, signal_791,
         signal_1583, signal_854, signal_1434, signal_790, signal_1585,
         signal_853, signal_1433, signal_789, signal_1587, signal_852,
         signal_1432, signal_788, signal_1589, signal_851, signal_1431,
         signal_787, signal_1591, signal_850, signal_1430, signal_786,
         signal_1593, signal_849, signal_1429, signal_785, signal_1595,
         signal_848, signal_1428, signal_784, signal_1597, signal_847,
         signal_1427, signal_783, signal_1599, signal_846, signal_1426,
         signal_782, signal_1601, signal_845, signal_1425, signal_781,
         signal_1603, signal_844, signal_1424, signal_780, signal_1605,
         signal_843, signal_1423, signal_779, signal_1607, signal_842,
         signal_1422, signal_778, signal_1609, signal_841, signal_1421,
         signal_777, signal_1611, signal_840, signal_1420, signal_776, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, cell_1001_n7,
         cell_1001_n6, cell_1001_n5, cell_1001_n3, cell_1001_n2, cell_1001_n1,
         cell_1001_LatchedEnable, cell_1001_N5, cell_1001_ShiftRegister_3_,
         cell_1000_n176, cell_1000_n175, cell_1000_n174, cell_1000_n173,
         cell_1000_n172, cell_1000_n171, cell_1000_n170, cell_1000_n169,
         cell_1000_n168, cell_1000_n167, cell_1000_n166, cell_1000_n165,
         cell_1000_n164, cell_1000_n163, cell_1000_n162, cell_1000_n161,
         cell_1000_n160, cell_1000_n159, cell_1000_n158, cell_1000_n157,
         cell_1000_n156, cell_1000_n155, cell_1000_n154, cell_1000_n153,
         cell_1000_n152, cell_1000_n151, cell_1000_n150, cell_1000_n149,
         cell_1000_n148, cell_1000_n147, cell_1000_n146, cell_1000_n145,
         cell_1000_n144, cell_1000_n143, cell_1000_n142, cell_1000_n141,
         cell_1000_n140, cell_1000_n139, cell_1000_n138, cell_1000_n137,
         cell_1000_n136, cell_1000_n135, cell_1000_n134, cell_1000_n133,
         cell_1000_n132, cell_1000_n131, cell_1000_n130, cell_1000_n129,
         cell_1000_n128, cell_1000_n127, cell_1000_n126, cell_1000_n125,
         cell_1000_n124, cell_1000_n123, cell_1000_n122, cell_1000_n121,
         cell_1000_n120, cell_1000_n119, cell_1000_n118, cell_1000_n117,
         cell_1000_n116, cell_1000_n115, cell_1000_n114, cell_1000_n113,
         cell_1000_n112, cell_1000_n111, cell_1000_n110, cell_1000_n109,
         cell_1000_n108, cell_1000_n107, cell_1000_n106, cell_1000_n105,
         cell_1000_n104, cell_1000_n103, cell_1000_n102, cell_1000_n101,
         cell_1000_n100, cell_1000_n99, cell_1000_n98, cell_1000_n97,
         cell_1000_n96, cell_1000_n95, cell_1000_n94, cell_1000_n93,
         cell_1000_n92, cell_1000_n91, cell_1000_n90, cell_1000_n89,
         cell_1000_n88, cell_1000_n87, cell_1000_n86, cell_1000_n85,
         cell_1000_n84, cell_1000_n83, cell_1000_n82, cell_1000_n81,
         cell_1000_n80, cell_1000_n79, cell_1000_n78, cell_1000_n77,
         cell_1000_n76, cell_1000_n75, cell_1000_n74, cell_1000_n73,
         cell_1000_n72, cell_1000_n71, cell_1000_n70, cell_1000_n69,
         cell_1000_n68, cell_1000_n67, cell_1000_n66, cell_1000_n65,
         cell_1000_n64, cell_1000_n63, cell_1000_n62, cell_1000_n61,
         cell_1000_n60, cell_1000_n59, cell_1000_n58, cell_1000_n57,
         cell_1000_n56, cell_1000_n55, cell_1000_n54, cell_1000_n53,
         cell_1000_n52, cell_1000_n51, cell_1000_n50, cell_1000_n49,
         cell_1000_n48, cell_1000_n47, cell_1000_n46, cell_1000_n45,
         cell_1000_n44, cell_1000_n43, cell_1000_n42, cell_1000_n41,
         cell_1000_n40, cell_1000_n39, cell_1000_n38, cell_1000_n37,
         cell_1000_n36, cell_1000_n35, cell_1000_n34, cell_1000_n33,
         cell_1000_n32, cell_1000_n31, cell_1000_n30, cell_1000_n29,
         cell_1000_n28, cell_1000_n27, cell_1000_n26, cell_1000_n25,
         cell_1000_n24, cell_1000_n23, cell_1000_n22, cell_1000_n21,
         cell_1000_n20, cell_1000_n19, cell_1000_n18, cell_1000_n17,
         cell_1000_n16, cell_1000_n15, cell_1000_n14, cell_1000_n13,
         cell_1000_n12, cell_1000_n11, cell_1000_n10, cell_1000_n9,
         cell_1000_n8, cell_1000_n7, cell_1000_n6, cell_1000_n5, cell_1000_n4,
         cell_1000_n3, cell_1000_n2, cell_1000_n1, cell_1000_g14_1_0_,
         cell_1000_g14_1_1_, cell_1000_g14_1_2_, cell_1000_g14_1_3_,
         cell_1000_g14_0_0_, cell_1000_g14_0_1_, cell_1000_g14_0_2_,
         cell_1000_g14_0_3_, cell_1000_g13_1_0_, cell_1000_g13_1_1_,
         cell_1000_g13_1_2_, cell_1000_g13_1_3_, cell_1000_g13_0_0_,
         cell_1000_g13_0_1_, cell_1000_g13_0_2_, cell_1000_g13_0_3_,
         cell_1000_g12_1_0_, cell_1000_g12_1_1_, cell_1000_g12_1_2_,
         cell_1000_g12_1_3_, cell_1000_g12_0_0_, cell_1000_g12_0_1_,
         cell_1000_g12_0_2_, cell_1000_g12_0_3_, cell_1000_g11_1_0_,
         cell_1000_g11_1_1_, cell_1000_g11_1_2_, cell_1000_g11_1_3_,
         cell_1000_g11_0_0_, cell_1000_g11_0_1_, cell_1000_g11_0_2_,
         cell_1000_g11_0_3_, cell_1000_g10_1_0_, cell_1000_g10_1_1_,
         cell_1000_g10_1_2_, cell_1000_g10_1_3_, cell_1000_g10_0_0_,
         cell_1000_g10_0_1_, cell_1000_g10_0_2_, cell_1000_g10_0_3_,
         cell_1000_g9_1_0_, cell_1000_g9_1_1_, cell_1000_g9_1_2_,
         cell_1000_g9_1_3_, cell_1000_g9_0_0_, cell_1000_g9_0_1_,
         cell_1000_g9_0_2_, cell_1000_g9_0_3_, cell_1000_g8_1_0_,
         cell_1000_g8_1_1_, cell_1000_g8_1_2_, cell_1000_g8_1_3_,
         cell_1000_g8_0_0_, cell_1000_g8_0_1_, cell_1000_g8_0_2_,
         cell_1000_g8_0_3_, cell_1000_g7_1_0_, cell_1000_g7_1_1_,
         cell_1000_g7_1_2_, cell_1000_g7_1_3_, cell_1000_g7_0_0_,
         cell_1000_g7_0_1_, cell_1000_g7_0_2_, cell_1000_g7_0_3_,
         cell_1000_g6_1_0_, cell_1000_g6_1_1_, cell_1000_g6_1_2_,
         cell_1000_g6_1_3_, cell_1000_g6_0_0_, cell_1000_g6_0_1_,
         cell_1000_g6_0_2_, cell_1000_g6_0_3_, cell_1000_g5_1_0_,
         cell_1000_g5_1_1_, cell_1000_g5_1_2_, cell_1000_g5_1_3_,
         cell_1000_g5_0_0_, cell_1000_g5_0_1_, cell_1000_g5_0_2_,
         cell_1000_g5_0_3_, cell_1000_g4_1_0_, cell_1000_g4_1_1_,
         cell_1000_g4_1_2_, cell_1000_g4_1_3_, cell_1000_g4_0_0_,
         cell_1000_g4_0_1_, cell_1000_g4_0_2_, cell_1000_g4_0_3_,
         cell_1000_g3_1_0_, cell_1000_g3_1_1_, cell_1000_g3_1_2_,
         cell_1000_g3_1_3_, cell_1000_g3_0_0_, cell_1000_g3_0_1_,
         cell_1000_g3_0_2_, cell_1000_g3_0_3_, cell_1000_g2_1_0_,
         cell_1000_g2_1_1_, cell_1000_g2_1_2_, cell_1000_g2_1_3_,
         cell_1000_g2_0_0_, cell_1000_g2_0_1_, cell_1000_g2_0_2_,
         cell_1000_g2_0_3_, cell_1000_g1_1_0_, cell_1000_g1_1_1_,
         cell_1000_g1_1_2_, cell_1000_g1_1_3_, cell_1000_g1_0_0_,
         cell_1000_g1_0_1_, cell_1000_g1_0_2_, cell_1000_g1_0_3_,
         cell_1000_g0_1_0_, cell_1000_g0_1_1_, cell_1000_g0_1_2_,
         cell_1000_g0_1_3_, cell_1000_g0_0_0_, cell_1000_g0_0_1_,
         cell_1000_g0_0_2_, cell_1000_g0_0_3_,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n379,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n378,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n377,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n376,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n375,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n373,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n372,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n368,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n367,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n366,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n365,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n363,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n360,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n358,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n225,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n224,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n223,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n222,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n221,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n220,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n219,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n218,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n217,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n216,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n215,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n213,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n212,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n211,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n210,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n180,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n179,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n178,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n177,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n176,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n15,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n14,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n13,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n12,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n68,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n67,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n379,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n378,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n377,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n376,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n375,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n373,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n372,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n368,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n367,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n366,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n365,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n363,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n360,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n358,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n225,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n224,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n223,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n222,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n221,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n220,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n219,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n218,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n217,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n216,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n215,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n213,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n212,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n211,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n210,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n180,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n179,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n178,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n177,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n176,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n15,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n14,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n13,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n12,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n379,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n378,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n377,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n376,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n375,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n373,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n372,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n368,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n367,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n366,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n365,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n363,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n360,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n358,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n225,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n224,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n223,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n222,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n221,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n220,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n219,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n218,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n217,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n216,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n215,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n213,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n212,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n211,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n210,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n180,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n179,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n178,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n177,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n176,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n15,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n14,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n13,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n12,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n379,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n378,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n377,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n376,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n375,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n373,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n372,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n368,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n367,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n366,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n365,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n363,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n360,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n358,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n225,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n224,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n223,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n222,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n221,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n220,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n219,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n218,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n217,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n216,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n215,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n213,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n212,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n211,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n210,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n180,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n179,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n178,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n177,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n176,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n15,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n14,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n13,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n12,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n379,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n378,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n377,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n376,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n375,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n373,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n372,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n368,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n367,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n366,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n365,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n363,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n360,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n358,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n225,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n224,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n223,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n222,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n221,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n220,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n219,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n218,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n217,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n216,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n215,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n213,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n212,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n211,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n210,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n180,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n179,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n178,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n177,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n176,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n15,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n14,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n13,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n12,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n379,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n378,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n377,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n376,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n375,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n373,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n372,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n368,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n367,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n366,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n365,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n363,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n360,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n358,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n225,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n224,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n223,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n222,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n221,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n220,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n219,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n218,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n217,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n216,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n215,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n213,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n212,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n211,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n210,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n180,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n179,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n178,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n177,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n176,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n15,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n14,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n13,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n12,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n379,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n378,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n377,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n376,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n375,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n373,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n372,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n368,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n367,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n366,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n365,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n363,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n360,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n358,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n225,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n224,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n223,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n222,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n221,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n220,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n219,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n218,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n217,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n216,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n215,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n213,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n212,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n211,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n210,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n180,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n179,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n178,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n177,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n176,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n15,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n14,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n13,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n12,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n379,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n378,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n377,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n376,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n375,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n373,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n372,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n368,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n367,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n366,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n365,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n363,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n360,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n358,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n225,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n224,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n223,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n222,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n221,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n220,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n219,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n218,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n217,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n216,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n215,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n213,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n212,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n211,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n210,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n180,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n179,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n178,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n177,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n176,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n15,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n14,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n13,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n12,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n379,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n378,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n377,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n376,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n375,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n373,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n372,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n368,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n367,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n366,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n365,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n363,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n360,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n358,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n225,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n224,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n223,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n222,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n221,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n220,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n219,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n218,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n217,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n216,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n215,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n213,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n212,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n211,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n210,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n180,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n179,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n178,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n177,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n176,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n15,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n14,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n13,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n12,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n379,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n378,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n377,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n376,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n375,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n373,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n372,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n368,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n367,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n366,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n365,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n363,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n360,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n358,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n225,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n224,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n223,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n222,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n221,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n220,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n219,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n218,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n217,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n216,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n215,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n213,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n212,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n211,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n210,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n180,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n179,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n178,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n177,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n176,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n15,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n14,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n13,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n12,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n379,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n378,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n377,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n376,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n375,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n373,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n372,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n368,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n367,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n366,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n365,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n363,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n360,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n358,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n225,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n224,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n223,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n222,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n221,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n220,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n219,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n218,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n217,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n216,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n215,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n213,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n212,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n211,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n210,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n180,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n179,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n178,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n177,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n176,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n15,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n14,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n13,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n12,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n379,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n378,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n377,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n376,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n375,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n373,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n372,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n368,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n367,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n366,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n365,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n363,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n360,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n358,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n225,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n224,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n223,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n222,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n221,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n220,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n219,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n218,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n217,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n216,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n215,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n213,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n212,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n211,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n210,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n180,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n179,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n178,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n177,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n176,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n15,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n14,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n13,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n12,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n379,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n378,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n377,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n376,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n375,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n373,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n372,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n368,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n367,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n366,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n365,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n363,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n360,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n358,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n225,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n224,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n223,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n222,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n221,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n220,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n219,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n218,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n217,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n216,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n215,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n213,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n212,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n211,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n210,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n180,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n179,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n178,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n177,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n176,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n15,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n14,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n13,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n12,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n379,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n378,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n377,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n376,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n375,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n373,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n372,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n368,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n367,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n366,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n365,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n363,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n360,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n358,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n225,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n224,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n223,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n222,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n221,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n220,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n219,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n218,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n217,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n216,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n215,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n213,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n212,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n211,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n210,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n180,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n179,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n178,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n177,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n176,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n15,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n14,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n13,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n12,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n379,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n378,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n377,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n376,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n375,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n373,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n372,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n368,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n367,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n366,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n365,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n363,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n360,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n358,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n225,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n224,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n223,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n222,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n221,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n220,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n219,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n218,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n217,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n216,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n215,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n213,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n212,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n211,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n210,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n180,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n179,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n178,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n177,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n176,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n15,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n14,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n13,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n12,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_15_value,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n379,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n378,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n377,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n376,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n375,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n373,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n372,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n368,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n367,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n366,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n365,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n363,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n360,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n358,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n225,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n224,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n223,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n222,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n221,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n220,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n219,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n218,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n217,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n216,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n215,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n213,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n212,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n211,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n210,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n180,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n179,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n178,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n177,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n176,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n15,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n14,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n13,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n12,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n232,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n231,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n230,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n229,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n228,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n227,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n226,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n225,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n224,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n223,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n222,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n221,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n220,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n219,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n218,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n217,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n216,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n215,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n214,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n213,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n212,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n211,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n210,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n209,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n208,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n207,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n206,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n205,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n204,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n203,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n202,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n201,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_0_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_1_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_2_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_3_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_4_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_5_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_6_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_7_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_8_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_9_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_10_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_11_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_12_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_13_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_14_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_15_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_0_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_1_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_2_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_3_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_4_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_5_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_6_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_7_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_8_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_9_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_10_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_11_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_12_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_13_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_14_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_15_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_0_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_1_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_2_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_3_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_4_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_5_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_6_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_7_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_8_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_9_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_10_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_11_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_12_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_13_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_14_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_15_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_0_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_1_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_2_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_3_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_4_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_5_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_6_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_7_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_8_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_9_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_10_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_11_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_12_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_13_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_14_value,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_15_value;
  wire   [3:0] cell_1000_g15_1;
  wire   [3:0] cell_1000_g15_0;
  wire   [3:0] cell_1000_GHPC_Gadget_0_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_0_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_0_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_1_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_1_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_1_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_2_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_2_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_2_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_3_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_3_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_3_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_4_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_4_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_4_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_5_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_5_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_5_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_6_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_6_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_6_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_7_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_7_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_7_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_8_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_8_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_8_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_9_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_9_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_9_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_10_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_10_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_10_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_11_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_11_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_11_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_12_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_12_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_12_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_13_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_13_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_13_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_14_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_14_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_14_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_15_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_15_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_15_inst_in1_reg;
  wire   [46:0] cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1;
  wire   [63:0] cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg;

  DFF_X1 cell_968 ( .D(signal_1030), .CK(signal_1676), .Q(signal_939), .QN(n31) );
  DFF_X1 cell_970 ( .D(signal_1031), .CK(signal_1676), .Q(signal_940), .QN(n29) );
  DFF_X1 cell_972 ( .D(signal_1032), .CK(signal_1676), .Q(signal_1025), .QN()
         );
  DFF_X1 cell_974 ( .D(signal_1033), .CK(signal_1676), .Q(signal_1026), .QN()
         );
  DFF_X1 cell_976 ( .D(signal_1034), .CK(signal_1676), .Q(signal_943), .QN(n30) );
  DFF_X1 cell_978 ( .D(signal_1035), .CK(signal_1676), .Q(signal_1028), .QN()
         );
  NOR4_X1 U40 ( .A1(signal_1026), .A2(signal_943), .A3(signal_1025), .A4(n29), 
        .ZN(n28) );
  AND3_X1 U41 ( .A1(signal_1028), .A2(signal_939), .A3(n28), .ZN(done) );
  INV_X1 U42 ( .A(rst), .ZN(n32) );
  AND2_X1 U43 ( .A1(n32), .A2(signal_1028), .ZN(signal_1034) );
  NOR3_X1 U44 ( .A1(signal_1025), .A2(signal_1026), .A3(n30), .ZN(n36) );
  NAND3_X1 U45 ( .A1(signal_939), .A2(n36), .A3(signal_1034), .ZN(n33) );
  OAI21_X1 U46 ( .B1(rst), .B2(n29), .A(n33), .ZN(signal_1030) );
  AND2_X1 U47 ( .A1(n32), .A2(signal_1025), .ZN(signal_1031) );
  AND2_X1 U48 ( .A1(n32), .A2(signal_1026), .ZN(signal_1032) );
  NAND3_X1 U49 ( .A1(signal_939), .A2(signal_1028), .A3(n29), .ZN(n34) );
  AOI211_X1 U50 ( .C1(n32), .C2(n34), .A(signal_1032), .B(signal_1031), .ZN(
        n35) );
  NOR2_X1 U51 ( .A1(n35), .A2(n30), .ZN(signal_1033) );
  AOI21_X1 U52 ( .B1(n36), .B2(signal_1028), .A(signal_940), .ZN(n37) );
  OAI221_X1 U53 ( .B1(signal_939), .B2(signal_940), .C1(n31), .C2(n37), .A(n32), .ZN(signal_1035) );
  MUX2_X1 cell_769_Ins_0_U1 ( .A(signal_1163), .B(Key_s0[0]), .S(rst), .Z(
        signal_1099) );
  MUX2_X1 cell_769_Ins_1_U1 ( .A(signal_1164), .B(Key_s1[0]), .S(rst), .Z(
        signal_1166) );
  MUX2_X1 cell_770_Ins_0_U1 ( .A(signal_1162), .B(Key_s0[1]), .S(rst), .Z(
        signal_1098) );
  MUX2_X1 cell_770_Ins_1_U1 ( .A(signal_1167), .B(Key_s1[1]), .S(rst), .Z(
        signal_1169) );
  MUX2_X1 cell_771_Ins_0_U1 ( .A(signal_1161), .B(Key_s0[2]), .S(rst), .Z(
        signal_1097) );
  MUX2_X1 cell_771_Ins_1_U1 ( .A(signal_1170), .B(Key_s1[2]), .S(rst), .Z(
        signal_1172) );
  MUX2_X1 cell_772_Ins_0_U1 ( .A(signal_1160), .B(Key_s0[3]), .S(rst), .Z(
        signal_1096) );
  MUX2_X1 cell_772_Ins_1_U1 ( .A(signal_1173), .B(Key_s1[3]), .S(rst), .Z(
        signal_1175) );
  MUX2_X1 cell_773_Ins_0_U1 ( .A(signal_1159), .B(Key_s0[4]), .S(rst), .Z(
        signal_1095) );
  MUX2_X1 cell_773_Ins_1_U1 ( .A(signal_1176), .B(Key_s1[4]), .S(rst), .Z(
        signal_1178) );
  MUX2_X1 cell_774_Ins_0_U1 ( .A(signal_1158), .B(Key_s0[5]), .S(rst), .Z(
        signal_1094) );
  MUX2_X1 cell_774_Ins_1_U1 ( .A(signal_1179), .B(Key_s1[5]), .S(rst), .Z(
        signal_1181) );
  MUX2_X1 cell_775_Ins_0_U1 ( .A(signal_1157), .B(Key_s0[6]), .S(rst), .Z(
        signal_1093) );
  MUX2_X1 cell_775_Ins_1_U1 ( .A(signal_1182), .B(Key_s1[6]), .S(rst), .Z(
        signal_1184) );
  MUX2_X1 cell_776_Ins_0_U1 ( .A(signal_1156), .B(Key_s0[7]), .S(rst), .Z(
        signal_1092) );
  MUX2_X1 cell_776_Ins_1_U1 ( .A(signal_1185), .B(Key_s1[7]), .S(rst), .Z(
        signal_1187) );
  MUX2_X1 cell_777_Ins_0_U1 ( .A(signal_1155), .B(Key_s0[8]), .S(rst), .Z(
        signal_1091) );
  MUX2_X1 cell_777_Ins_1_U1 ( .A(signal_1188), .B(Key_s1[8]), .S(rst), .Z(
        signal_1190) );
  MUX2_X1 cell_778_Ins_0_U1 ( .A(signal_1154), .B(Key_s0[9]), .S(rst), .Z(
        signal_1090) );
  MUX2_X1 cell_778_Ins_1_U1 ( .A(signal_1191), .B(Key_s1[9]), .S(rst), .Z(
        signal_1193) );
  MUX2_X1 cell_779_Ins_0_U1 ( .A(signal_1153), .B(Key_s0[10]), .S(rst), .Z(
        signal_1089) );
  MUX2_X1 cell_779_Ins_1_U1 ( .A(signal_1194), .B(Key_s1[10]), .S(rst), .Z(
        signal_1196) );
  MUX2_X1 cell_780_Ins_0_U1 ( .A(signal_1152), .B(Key_s0[11]), .S(rst), .Z(
        signal_1088) );
  MUX2_X1 cell_780_Ins_1_U1 ( .A(signal_1197), .B(Key_s1[11]), .S(rst), .Z(
        signal_1199) );
  MUX2_X1 cell_781_Ins_0_U1 ( .A(signal_1151), .B(Key_s0[12]), .S(rst), .Z(
        signal_1087) );
  MUX2_X1 cell_781_Ins_1_U1 ( .A(signal_1200), .B(Key_s1[12]), .S(rst), .Z(
        signal_1202) );
  MUX2_X1 cell_782_Ins_0_U1 ( .A(signal_1150), .B(Key_s0[13]), .S(rst), .Z(
        signal_1086) );
  MUX2_X1 cell_782_Ins_1_U1 ( .A(signal_1203), .B(Key_s1[13]), .S(rst), .Z(
        signal_1205) );
  MUX2_X1 cell_783_Ins_0_U1 ( .A(signal_1149), .B(Key_s0[14]), .S(rst), .Z(
        signal_1085) );
  MUX2_X1 cell_783_Ins_1_U1 ( .A(signal_1206), .B(Key_s1[14]), .S(rst), .Z(
        signal_1208) );
  MUX2_X1 cell_784_Ins_0_U1 ( .A(signal_1148), .B(Key_s0[15]), .S(rst), .Z(
        signal_1084) );
  MUX2_X1 cell_784_Ins_1_U1 ( .A(signal_1209), .B(Key_s1[15]), .S(rst), .Z(
        signal_1211) );
  MUX2_X1 cell_785_Ins_0_U1 ( .A(signal_1147), .B(Key_s0[16]), .S(rst), .Z(
        signal_1083) );
  MUX2_X1 cell_785_Ins_1_U1 ( .A(signal_1212), .B(Key_s1[16]), .S(rst), .Z(
        signal_1214) );
  MUX2_X1 cell_786_Ins_0_U1 ( .A(signal_1146), .B(Key_s0[17]), .S(rst), .Z(
        signal_1082) );
  MUX2_X1 cell_786_Ins_1_U1 ( .A(signal_1215), .B(Key_s1[17]), .S(rst), .Z(
        signal_1217) );
  MUX2_X1 cell_787_Ins_0_U1 ( .A(signal_1145), .B(Key_s0[18]), .S(rst), .Z(
        signal_1081) );
  MUX2_X1 cell_787_Ins_1_U1 ( .A(signal_1218), .B(Key_s1[18]), .S(rst), .Z(
        signal_1220) );
  MUX2_X1 cell_788_Ins_0_U1 ( .A(signal_1144), .B(Key_s0[19]), .S(rst), .Z(
        signal_1080) );
  MUX2_X1 cell_788_Ins_1_U1 ( .A(signal_1221), .B(Key_s1[19]), .S(rst), .Z(
        signal_1223) );
  MUX2_X1 cell_789_Ins_0_U1 ( .A(signal_1143), .B(Key_s0[20]), .S(rst), .Z(
        signal_1079) );
  MUX2_X1 cell_789_Ins_1_U1 ( .A(signal_1224), .B(Key_s1[20]), .S(rst), .Z(
        signal_1226) );
  MUX2_X1 cell_790_Ins_0_U1 ( .A(signal_1142), .B(Key_s0[21]), .S(rst), .Z(
        signal_1078) );
  MUX2_X1 cell_790_Ins_1_U1 ( .A(signal_1227), .B(Key_s1[21]), .S(rst), .Z(
        signal_1229) );
  MUX2_X1 cell_791_Ins_0_U1 ( .A(signal_1141), .B(Key_s0[22]), .S(rst), .Z(
        signal_1077) );
  MUX2_X1 cell_791_Ins_1_U1 ( .A(signal_1230), .B(Key_s1[22]), .S(rst), .Z(
        signal_1232) );
  MUX2_X1 cell_792_Ins_0_U1 ( .A(signal_1140), .B(Key_s0[23]), .S(rst), .Z(
        signal_1076) );
  MUX2_X1 cell_792_Ins_1_U1 ( .A(signal_1233), .B(Key_s1[23]), .S(rst), .Z(
        signal_1235) );
  MUX2_X1 cell_793_Ins_0_U1 ( .A(signal_1139), .B(Key_s0[24]), .S(rst), .Z(
        signal_1075) );
  MUX2_X1 cell_793_Ins_1_U1 ( .A(signal_1236), .B(Key_s1[24]), .S(rst), .Z(
        signal_1238) );
  MUX2_X1 cell_794_Ins_0_U1 ( .A(signal_1138), .B(Key_s0[25]), .S(rst), .Z(
        signal_1074) );
  MUX2_X1 cell_794_Ins_1_U1 ( .A(signal_1239), .B(Key_s1[25]), .S(rst), .Z(
        signal_1241) );
  MUX2_X1 cell_795_Ins_0_U1 ( .A(signal_1137), .B(Key_s0[26]), .S(rst), .Z(
        signal_1073) );
  MUX2_X1 cell_795_Ins_1_U1 ( .A(signal_1242), .B(Key_s1[26]), .S(rst), .Z(
        signal_1244) );
  MUX2_X1 cell_796_Ins_0_U1 ( .A(signal_1136), .B(Key_s0[27]), .S(rst), .Z(
        signal_1072) );
  MUX2_X1 cell_796_Ins_1_U1 ( .A(signal_1245), .B(Key_s1[27]), .S(rst), .Z(
        signal_1247) );
  MUX2_X1 cell_797_Ins_0_U1 ( .A(signal_1135), .B(Key_s0[28]), .S(rst), .Z(
        signal_1071) );
  MUX2_X1 cell_797_Ins_1_U1 ( .A(signal_1248), .B(Key_s1[28]), .S(rst), .Z(
        signal_1250) );
  MUX2_X1 cell_798_Ins_0_U1 ( .A(signal_1134), .B(Key_s0[29]), .S(rst), .Z(
        signal_1070) );
  MUX2_X1 cell_798_Ins_1_U1 ( .A(signal_1251), .B(Key_s1[29]), .S(rst), .Z(
        signal_1253) );
  MUX2_X1 cell_799_Ins_0_U1 ( .A(signal_1133), .B(Key_s0[30]), .S(rst), .Z(
        signal_1069) );
  MUX2_X1 cell_799_Ins_1_U1 ( .A(signal_1254), .B(Key_s1[30]), .S(rst), .Z(
        signal_1256) );
  MUX2_X1 cell_800_Ins_0_U1 ( .A(signal_1132), .B(Key_s0[31]), .S(rst), .Z(
        signal_1068) );
  MUX2_X1 cell_800_Ins_1_U1 ( .A(signal_1257), .B(Key_s1[31]), .S(rst), .Z(
        signal_1259) );
  MUX2_X1 cell_801_Ins_0_U1 ( .A(signal_1131), .B(Key_s0[32]), .S(rst), .Z(
        signal_1067) );
  MUX2_X1 cell_801_Ins_1_U1 ( .A(signal_1260), .B(Key_s1[32]), .S(rst), .Z(
        signal_1262) );
  MUX2_X1 cell_802_Ins_0_U1 ( .A(signal_1130), .B(Key_s0[33]), .S(rst), .Z(
        signal_1066) );
  MUX2_X1 cell_802_Ins_1_U1 ( .A(signal_1263), .B(Key_s1[33]), .S(rst), .Z(
        signal_1265) );
  MUX2_X1 cell_803_Ins_0_U1 ( .A(signal_1129), .B(Key_s0[34]), .S(rst), .Z(
        signal_1065) );
  MUX2_X1 cell_803_Ins_1_U1 ( .A(signal_1266), .B(Key_s1[34]), .S(rst), .Z(
        signal_1268) );
  MUX2_X1 cell_804_Ins_0_U1 ( .A(signal_1128), .B(Key_s0[35]), .S(rst), .Z(
        signal_1064) );
  MUX2_X1 cell_804_Ins_1_U1 ( .A(signal_1269), .B(Key_s1[35]), .S(rst), .Z(
        signal_1271) );
  MUX2_X1 cell_805_Ins_0_U1 ( .A(signal_1127), .B(Key_s0[36]), .S(rst), .Z(
        signal_1063) );
  MUX2_X1 cell_805_Ins_1_U1 ( .A(signal_1272), .B(Key_s1[36]), .S(rst), .Z(
        signal_1274) );
  MUX2_X1 cell_806_Ins_0_U1 ( .A(signal_1126), .B(Key_s0[37]), .S(rst), .Z(
        signal_1062) );
  MUX2_X1 cell_806_Ins_1_U1 ( .A(signal_1275), .B(Key_s1[37]), .S(rst), .Z(
        signal_1277) );
  MUX2_X1 cell_807_Ins_0_U1 ( .A(signal_1125), .B(Key_s0[38]), .S(rst), .Z(
        signal_1061) );
  MUX2_X1 cell_807_Ins_1_U1 ( .A(signal_1278), .B(Key_s1[38]), .S(rst), .Z(
        signal_1280) );
  MUX2_X1 cell_808_Ins_0_U1 ( .A(signal_1124), .B(Key_s0[39]), .S(rst), .Z(
        signal_1060) );
  MUX2_X1 cell_808_Ins_1_U1 ( .A(signal_1281), .B(Key_s1[39]), .S(rst), .Z(
        signal_1283) );
  MUX2_X1 cell_809_Ins_0_U1 ( .A(signal_1123), .B(Key_s0[40]), .S(rst), .Z(
        signal_1059) );
  MUX2_X1 cell_809_Ins_1_U1 ( .A(signal_1284), .B(Key_s1[40]), .S(rst), .Z(
        signal_1286) );
  MUX2_X1 cell_810_Ins_0_U1 ( .A(signal_1122), .B(Key_s0[41]), .S(rst), .Z(
        signal_1058) );
  MUX2_X1 cell_810_Ins_1_U1 ( .A(signal_1287), .B(Key_s1[41]), .S(rst), .Z(
        signal_1289) );
  MUX2_X1 cell_811_Ins_0_U1 ( .A(signal_1121), .B(Key_s0[42]), .S(rst), .Z(
        signal_1057) );
  MUX2_X1 cell_811_Ins_1_U1 ( .A(signal_1290), .B(Key_s1[42]), .S(rst), .Z(
        signal_1292) );
  MUX2_X1 cell_812_Ins_0_U1 ( .A(signal_1120), .B(Key_s0[43]), .S(rst), .Z(
        signal_1056) );
  MUX2_X1 cell_812_Ins_1_U1 ( .A(signal_1293), .B(Key_s1[43]), .S(rst), .Z(
        signal_1295) );
  MUX2_X1 cell_813_Ins_0_U1 ( .A(signal_1119), .B(Key_s0[44]), .S(rst), .Z(
        signal_1055) );
  MUX2_X1 cell_813_Ins_1_U1 ( .A(signal_1296), .B(Key_s1[44]), .S(rst), .Z(
        signal_1298) );
  MUX2_X1 cell_814_Ins_0_U1 ( .A(signal_1118), .B(Key_s0[45]), .S(rst), .Z(
        signal_1054) );
  MUX2_X1 cell_814_Ins_1_U1 ( .A(signal_1299), .B(Key_s1[45]), .S(rst), .Z(
        signal_1301) );
  MUX2_X1 cell_815_Ins_0_U1 ( .A(signal_1117), .B(Key_s0[46]), .S(rst), .Z(
        signal_1053) );
  MUX2_X1 cell_815_Ins_1_U1 ( .A(signal_1302), .B(Key_s1[46]), .S(rst), .Z(
        signal_1304) );
  MUX2_X1 cell_816_Ins_0_U1 ( .A(signal_1116), .B(Key_s0[47]), .S(rst), .Z(
        signal_1052) );
  MUX2_X1 cell_816_Ins_1_U1 ( .A(signal_1305), .B(Key_s1[47]), .S(rst), .Z(
        signal_1307) );
  MUX2_X1 cell_817_Ins_0_U1 ( .A(signal_1115), .B(Key_s0[48]), .S(rst), .Z(
        signal_1051) );
  MUX2_X1 cell_817_Ins_1_U1 ( .A(signal_1308), .B(Key_s1[48]), .S(rst), .Z(
        signal_1310) );
  MUX2_X1 cell_818_Ins_0_U1 ( .A(signal_1114), .B(Key_s0[49]), .S(rst), .Z(
        signal_1050) );
  MUX2_X1 cell_818_Ins_1_U1 ( .A(signal_1311), .B(Key_s1[49]), .S(rst), .Z(
        signal_1313) );
  MUX2_X1 cell_819_Ins_0_U1 ( .A(signal_1113), .B(Key_s0[50]), .S(rst), .Z(
        signal_1049) );
  MUX2_X1 cell_819_Ins_1_U1 ( .A(signal_1314), .B(Key_s1[50]), .S(rst), .Z(
        signal_1316) );
  MUX2_X1 cell_820_Ins_0_U1 ( .A(signal_1112), .B(Key_s0[51]), .S(rst), .Z(
        signal_1048) );
  MUX2_X1 cell_820_Ins_1_U1 ( .A(signal_1317), .B(Key_s1[51]), .S(rst), .Z(
        signal_1319) );
  MUX2_X1 cell_821_Ins_0_U1 ( .A(signal_1111), .B(Key_s0[52]), .S(rst), .Z(
        signal_1047) );
  MUX2_X1 cell_821_Ins_1_U1 ( .A(signal_1320), .B(Key_s1[52]), .S(rst), .Z(
        signal_1322) );
  MUX2_X1 cell_822_Ins_0_U1 ( .A(signal_1110), .B(Key_s0[53]), .S(rst), .Z(
        signal_1046) );
  MUX2_X1 cell_822_Ins_1_U1 ( .A(signal_1323), .B(Key_s1[53]), .S(rst), .Z(
        signal_1325) );
  MUX2_X1 cell_823_Ins_0_U1 ( .A(signal_1109), .B(Key_s0[54]), .S(rst), .Z(
        signal_1045) );
  MUX2_X1 cell_823_Ins_1_U1 ( .A(signal_1326), .B(Key_s1[54]), .S(rst), .Z(
        signal_1328) );
  MUX2_X1 cell_824_Ins_0_U1 ( .A(signal_1108), .B(Key_s0[55]), .S(rst), .Z(
        signal_1044) );
  MUX2_X1 cell_824_Ins_1_U1 ( .A(signal_1329), .B(Key_s1[55]), .S(rst), .Z(
        signal_1331) );
  MUX2_X1 cell_825_Ins_0_U1 ( .A(signal_1107), .B(Key_s0[56]), .S(rst), .Z(
        signal_1043) );
  MUX2_X1 cell_825_Ins_1_U1 ( .A(signal_1332), .B(Key_s1[56]), .S(rst), .Z(
        signal_1334) );
  MUX2_X1 cell_826_Ins_0_U1 ( .A(signal_1106), .B(Key_s0[57]), .S(rst), .Z(
        signal_1042) );
  MUX2_X1 cell_826_Ins_1_U1 ( .A(signal_1335), .B(Key_s1[57]), .S(rst), .Z(
        signal_1337) );
  MUX2_X1 cell_827_Ins_0_U1 ( .A(signal_1105), .B(Key_s0[58]), .S(rst), .Z(
        signal_1041) );
  MUX2_X1 cell_827_Ins_1_U1 ( .A(signal_1338), .B(Key_s1[58]), .S(rst), .Z(
        signal_1340) );
  MUX2_X1 cell_828_Ins_0_U1 ( .A(signal_1104), .B(Key_s0[59]), .S(rst), .Z(
        signal_1040) );
  MUX2_X1 cell_828_Ins_1_U1 ( .A(signal_1341), .B(Key_s1[59]), .S(rst), .Z(
        signal_1343) );
  MUX2_X1 cell_829_Ins_0_U1 ( .A(signal_1103), .B(Key_s0[60]), .S(rst), .Z(
        signal_1039) );
  MUX2_X1 cell_829_Ins_1_U1 ( .A(signal_1344), .B(Key_s1[60]), .S(rst), .Z(
        signal_1346) );
  MUX2_X1 cell_830_Ins_0_U1 ( .A(signal_1102), .B(Key_s0[61]), .S(rst), .Z(
        signal_1038) );
  MUX2_X1 cell_830_Ins_1_U1 ( .A(signal_1347), .B(Key_s1[61]), .S(rst), .Z(
        signal_1349) );
  MUX2_X1 cell_831_Ins_0_U1 ( .A(signal_1101), .B(Key_s0[62]), .S(rst), .Z(
        signal_1037) );
  MUX2_X1 cell_831_Ins_1_U1 ( .A(signal_1350), .B(Key_s1[62]), .S(rst), .Z(
        signal_1352) );
  MUX2_X1 cell_832_Ins_0_U1 ( .A(signal_1100), .B(Key_s0[63]), .S(rst), .Z(
        signal_1036) );
  MUX2_X1 cell_832_Ins_1_U1 ( .A(signal_1353), .B(Key_s1[63]), .S(rst), .Z(
        signal_1355) );
  NOR2_X1 cell_1001_U7 ( .A1(rst), .A2(cell_1001_n6), .ZN(cell_1001_n2) );
  NOR2_X1 cell_1001_U6 ( .A1(rst), .A2(cell_1001_n5), .ZN(cell_1001_n1) );
  NAND2_X1 cell_1001_U5 ( .A1(cell_1001_n3), .A2(cell_1001_n7), .ZN(
        cell_1001_N5) );
  AND2_X1 cell_1001_U4 ( .A1(cell_1001_LatchedEnable), .A2(clk), .ZN(
        signal_1676) );
  INV_X1 cell_1001_U3 ( .A(rst), .ZN(cell_1001_n7) );
  DFF_X1 cell_1001_ShiftRegister_reg_2_ ( .D(cell_1001_n1), .CK(clk), .Q(), 
        .QN(cell_1001_n6) );
  DFF_X1 cell_1001_ShiftRegister_reg_3_ ( .D(cell_1001_n2), .CK(clk), .Q(
        cell_1001_ShiftRegister_3_), .QN(cell_1001_n3) );
  DLL_X1 cell_1001_LatchedEnable_reg ( .D(cell_1001_N5), .GN(clk), .Q(
        cell_1001_LatchedEnable) );
  DLL_X1 cell_1001_Synch_reg ( .D(cell_1001_ShiftRegister_3_), .GN(clk), .Q(
        Synch) );
  DFF_X1 cell_1001_ShiftRegister_reg_1_ ( .D(cell_1001_N5), .CK(clk), .Q(), 
        .QN(cell_1001_n5) );
  MUX2_X1 cell_0_Ins_0_U1 ( .A(signal_839), .B(Plaintext_s0[0]), .S(rst), .Z(
        signal_903) );
  MUX2_X1 cell_0_Ins_1_U1 ( .A(signal_1483), .B(Plaintext_s1[0]), .S(rst), .Z(
        signal_1485) );
  MUX2_X1 cell_1_Ins_0_U1 ( .A(signal_838), .B(Plaintext_s0[1]), .S(rst), .Z(
        signal_902) );
  MUX2_X1 cell_1_Ins_1_U1 ( .A(signal_1482), .B(Plaintext_s1[1]), .S(rst), .Z(
        signal_1487) );
  MUX2_X1 cell_2_Ins_0_U1 ( .A(signal_837), .B(Plaintext_s0[2]), .S(rst), .Z(
        signal_901) );
  MUX2_X1 cell_2_Ins_1_U1 ( .A(signal_1481), .B(Plaintext_s1[2]), .S(rst), .Z(
        signal_1489) );
  MUX2_X1 cell_3_Ins_0_U1 ( .A(signal_836), .B(Plaintext_s0[3]), .S(rst), .Z(
        signal_900) );
  MUX2_X1 cell_3_Ins_1_U1 ( .A(signal_1480), .B(Plaintext_s1[3]), .S(rst), .Z(
        signal_1491) );
  MUX2_X1 cell_4_Ins_0_U1 ( .A(signal_835), .B(Plaintext_s0[4]), .S(rst), .Z(
        signal_899) );
  MUX2_X1 cell_4_Ins_1_U1 ( .A(signal_1479), .B(Plaintext_s1[4]), .S(rst), .Z(
        signal_1493) );
  MUX2_X1 cell_5_Ins_0_U1 ( .A(signal_834), .B(Plaintext_s0[5]), .S(rst), .Z(
        signal_898) );
  MUX2_X1 cell_5_Ins_1_U1 ( .A(signal_1478), .B(Plaintext_s1[5]), .S(rst), .Z(
        signal_1495) );
  MUX2_X1 cell_6_Ins_0_U1 ( .A(signal_833), .B(Plaintext_s0[6]), .S(rst), .Z(
        signal_897) );
  MUX2_X1 cell_6_Ins_1_U1 ( .A(signal_1477), .B(Plaintext_s1[6]), .S(rst), .Z(
        signal_1497) );
  MUX2_X1 cell_7_Ins_0_U1 ( .A(signal_832), .B(Plaintext_s0[7]), .S(rst), .Z(
        signal_896) );
  MUX2_X1 cell_7_Ins_1_U1 ( .A(signal_1476), .B(Plaintext_s1[7]), .S(rst), .Z(
        signal_1499) );
  MUX2_X1 cell_8_Ins_0_U1 ( .A(signal_831), .B(Plaintext_s0[8]), .S(rst), .Z(
        signal_895) );
  MUX2_X1 cell_8_Ins_1_U1 ( .A(signal_1475), .B(Plaintext_s1[8]), .S(rst), .Z(
        signal_1501) );
  MUX2_X1 cell_9_Ins_0_U1 ( .A(signal_830), .B(Plaintext_s0[9]), .S(rst), .Z(
        signal_894) );
  MUX2_X1 cell_9_Ins_1_U1 ( .A(signal_1474), .B(Plaintext_s1[9]), .S(rst), .Z(
        signal_1503) );
  MUX2_X1 cell_10_Ins_0_U1 ( .A(signal_829), .B(Plaintext_s0[10]), .S(rst), 
        .Z(signal_893) );
  MUX2_X1 cell_10_Ins_1_U1 ( .A(signal_1473), .B(Plaintext_s1[10]), .S(rst), 
        .Z(signal_1505) );
  MUX2_X1 cell_11_Ins_0_U1 ( .A(signal_828), .B(Plaintext_s0[11]), .S(rst), 
        .Z(signal_892) );
  MUX2_X1 cell_11_Ins_1_U1 ( .A(signal_1472), .B(Plaintext_s1[11]), .S(rst), 
        .Z(signal_1507) );
  MUX2_X1 cell_12_Ins_0_U1 ( .A(signal_827), .B(Plaintext_s0[12]), .S(rst), 
        .Z(signal_891) );
  MUX2_X1 cell_12_Ins_1_U1 ( .A(signal_1471), .B(Plaintext_s1[12]), .S(rst), 
        .Z(signal_1509) );
  MUX2_X1 cell_13_Ins_0_U1 ( .A(signal_826), .B(Plaintext_s0[13]), .S(rst), 
        .Z(signal_890) );
  MUX2_X1 cell_13_Ins_1_U1 ( .A(signal_1470), .B(Plaintext_s1[13]), .S(rst), 
        .Z(signal_1511) );
  MUX2_X1 cell_14_Ins_0_U1 ( .A(signal_825), .B(Plaintext_s0[14]), .S(rst), 
        .Z(signal_889) );
  MUX2_X1 cell_14_Ins_1_U1 ( .A(signal_1469), .B(Plaintext_s1[14]), .S(rst), 
        .Z(signal_1513) );
  MUX2_X1 cell_15_Ins_0_U1 ( .A(signal_824), .B(Plaintext_s0[15]), .S(rst), 
        .Z(signal_888) );
  MUX2_X1 cell_15_Ins_1_U1 ( .A(signal_1468), .B(Plaintext_s1[15]), .S(rst), 
        .Z(signal_1515) );
  MUX2_X1 cell_16_Ins_0_U1 ( .A(signal_823), .B(Plaintext_s0[16]), .S(rst), 
        .Z(signal_887) );
  MUX2_X1 cell_16_Ins_1_U1 ( .A(signal_1467), .B(Plaintext_s1[16]), .S(rst), 
        .Z(signal_1517) );
  MUX2_X1 cell_17_Ins_0_U1 ( .A(signal_822), .B(Plaintext_s0[17]), .S(rst), 
        .Z(signal_886) );
  MUX2_X1 cell_17_Ins_1_U1 ( .A(signal_1466), .B(Plaintext_s1[17]), .S(rst), 
        .Z(signal_1519) );
  MUX2_X1 cell_18_Ins_0_U1 ( .A(signal_821), .B(Plaintext_s0[18]), .S(rst), 
        .Z(signal_885) );
  MUX2_X1 cell_18_Ins_1_U1 ( .A(signal_1465), .B(Plaintext_s1[18]), .S(rst), 
        .Z(signal_1521) );
  MUX2_X1 cell_19_Ins_0_U1 ( .A(signal_820), .B(Plaintext_s0[19]), .S(rst), 
        .Z(signal_884) );
  MUX2_X1 cell_19_Ins_1_U1 ( .A(signal_1464), .B(Plaintext_s1[19]), .S(rst), 
        .Z(signal_1523) );
  MUX2_X1 cell_20_Ins_0_U1 ( .A(signal_819), .B(Plaintext_s0[20]), .S(rst), 
        .Z(signal_883) );
  MUX2_X1 cell_20_Ins_1_U1 ( .A(signal_1463), .B(Plaintext_s1[20]), .S(rst), 
        .Z(signal_1525) );
  MUX2_X1 cell_21_Ins_0_U1 ( .A(signal_818), .B(Plaintext_s0[21]), .S(rst), 
        .Z(signal_882) );
  MUX2_X1 cell_21_Ins_1_U1 ( .A(signal_1462), .B(Plaintext_s1[21]), .S(rst), 
        .Z(signal_1527) );
  MUX2_X1 cell_22_Ins_0_U1 ( .A(signal_817), .B(Plaintext_s0[22]), .S(rst), 
        .Z(signal_881) );
  MUX2_X1 cell_22_Ins_1_U1 ( .A(signal_1461), .B(Plaintext_s1[22]), .S(rst), 
        .Z(signal_1529) );
  MUX2_X1 cell_23_Ins_0_U1 ( .A(signal_816), .B(Plaintext_s0[23]), .S(rst), 
        .Z(signal_880) );
  MUX2_X1 cell_23_Ins_1_U1 ( .A(signal_1460), .B(Plaintext_s1[23]), .S(rst), 
        .Z(signal_1531) );
  MUX2_X1 cell_24_Ins_0_U1 ( .A(signal_815), .B(Plaintext_s0[24]), .S(rst), 
        .Z(signal_879) );
  MUX2_X1 cell_24_Ins_1_U1 ( .A(signal_1459), .B(Plaintext_s1[24]), .S(rst), 
        .Z(signal_1533) );
  MUX2_X1 cell_25_Ins_0_U1 ( .A(signal_814), .B(Plaintext_s0[25]), .S(rst), 
        .Z(signal_878) );
  MUX2_X1 cell_25_Ins_1_U1 ( .A(signal_1458), .B(Plaintext_s1[25]), .S(rst), 
        .Z(signal_1535) );
  MUX2_X1 cell_26_Ins_0_U1 ( .A(signal_813), .B(Plaintext_s0[26]), .S(rst), 
        .Z(signal_877) );
  MUX2_X1 cell_26_Ins_1_U1 ( .A(signal_1457), .B(Plaintext_s1[26]), .S(rst), 
        .Z(signal_1537) );
  MUX2_X1 cell_27_Ins_0_U1 ( .A(signal_812), .B(Plaintext_s0[27]), .S(rst), 
        .Z(signal_876) );
  MUX2_X1 cell_27_Ins_1_U1 ( .A(signal_1456), .B(Plaintext_s1[27]), .S(rst), 
        .Z(signal_1539) );
  MUX2_X1 cell_28_Ins_0_U1 ( .A(signal_811), .B(Plaintext_s0[28]), .S(rst), 
        .Z(signal_875) );
  MUX2_X1 cell_28_Ins_1_U1 ( .A(signal_1455), .B(Plaintext_s1[28]), .S(rst), 
        .Z(signal_1541) );
  MUX2_X1 cell_29_Ins_0_U1 ( .A(signal_810), .B(Plaintext_s0[29]), .S(rst), 
        .Z(signal_874) );
  MUX2_X1 cell_29_Ins_1_U1 ( .A(signal_1454), .B(Plaintext_s1[29]), .S(rst), 
        .Z(signal_1543) );
  MUX2_X1 cell_30_Ins_0_U1 ( .A(signal_809), .B(Plaintext_s0[30]), .S(rst), 
        .Z(signal_873) );
  MUX2_X1 cell_30_Ins_1_U1 ( .A(signal_1453), .B(Plaintext_s1[30]), .S(rst), 
        .Z(signal_1545) );
  MUX2_X1 cell_31_Ins_0_U1 ( .A(signal_808), .B(Plaintext_s0[31]), .S(rst), 
        .Z(signal_872) );
  MUX2_X1 cell_31_Ins_1_U1 ( .A(signal_1452), .B(Plaintext_s1[31]), .S(rst), 
        .Z(signal_1547) );
  MUX2_X1 cell_32_Ins_0_U1 ( .A(signal_807), .B(Plaintext_s0[32]), .S(rst), 
        .Z(signal_871) );
  MUX2_X1 cell_32_Ins_1_U1 ( .A(signal_1451), .B(Plaintext_s1[32]), .S(rst), 
        .Z(signal_1549) );
  MUX2_X1 cell_33_Ins_0_U1 ( .A(signal_806), .B(Plaintext_s0[33]), .S(rst), 
        .Z(signal_870) );
  MUX2_X1 cell_33_Ins_1_U1 ( .A(signal_1450), .B(Plaintext_s1[33]), .S(rst), 
        .Z(signal_1551) );
  MUX2_X1 cell_34_Ins_0_U1 ( .A(signal_805), .B(Plaintext_s0[34]), .S(rst), 
        .Z(signal_869) );
  MUX2_X1 cell_34_Ins_1_U1 ( .A(signal_1449), .B(Plaintext_s1[34]), .S(rst), 
        .Z(signal_1553) );
  MUX2_X1 cell_35_Ins_0_U1 ( .A(signal_804), .B(Plaintext_s0[35]), .S(rst), 
        .Z(signal_868) );
  MUX2_X1 cell_35_Ins_1_U1 ( .A(signal_1448), .B(Plaintext_s1[35]), .S(rst), 
        .Z(signal_1555) );
  MUX2_X1 cell_36_Ins_0_U1 ( .A(signal_803), .B(Plaintext_s0[36]), .S(rst), 
        .Z(signal_867) );
  MUX2_X1 cell_36_Ins_1_U1 ( .A(signal_1447), .B(Plaintext_s1[36]), .S(rst), 
        .Z(signal_1557) );
  MUX2_X1 cell_37_Ins_0_U1 ( .A(signal_802), .B(Plaintext_s0[37]), .S(rst), 
        .Z(signal_866) );
  MUX2_X1 cell_37_Ins_1_U1 ( .A(signal_1446), .B(Plaintext_s1[37]), .S(rst), 
        .Z(signal_1559) );
  MUX2_X1 cell_38_Ins_0_U1 ( .A(signal_801), .B(Plaintext_s0[38]), .S(rst), 
        .Z(signal_865) );
  MUX2_X1 cell_38_Ins_1_U1 ( .A(signal_1445), .B(Plaintext_s1[38]), .S(rst), 
        .Z(signal_1561) );
  MUX2_X1 cell_39_Ins_0_U1 ( .A(signal_800), .B(Plaintext_s0[39]), .S(rst), 
        .Z(signal_864) );
  MUX2_X1 cell_39_Ins_1_U1 ( .A(signal_1444), .B(Plaintext_s1[39]), .S(rst), 
        .Z(signal_1563) );
  MUX2_X1 cell_40_Ins_0_U1 ( .A(signal_799), .B(Plaintext_s0[40]), .S(rst), 
        .Z(signal_863) );
  MUX2_X1 cell_40_Ins_1_U1 ( .A(signal_1443), .B(Plaintext_s1[40]), .S(rst), 
        .Z(signal_1565) );
  MUX2_X1 cell_41_Ins_0_U1 ( .A(signal_798), .B(Plaintext_s0[41]), .S(rst), 
        .Z(signal_862) );
  MUX2_X1 cell_41_Ins_1_U1 ( .A(signal_1442), .B(Plaintext_s1[41]), .S(rst), 
        .Z(signal_1567) );
  MUX2_X1 cell_42_Ins_0_U1 ( .A(signal_797), .B(Plaintext_s0[42]), .S(rst), 
        .Z(signal_861) );
  MUX2_X1 cell_42_Ins_1_U1 ( .A(signal_1441), .B(Plaintext_s1[42]), .S(rst), 
        .Z(signal_1569) );
  MUX2_X1 cell_43_Ins_0_U1 ( .A(signal_796), .B(Plaintext_s0[43]), .S(rst), 
        .Z(signal_860) );
  MUX2_X1 cell_43_Ins_1_U1 ( .A(signal_1440), .B(Plaintext_s1[43]), .S(rst), 
        .Z(signal_1571) );
  MUX2_X1 cell_44_Ins_0_U1 ( .A(signal_795), .B(Plaintext_s0[44]), .S(rst), 
        .Z(signal_859) );
  MUX2_X1 cell_44_Ins_1_U1 ( .A(signal_1439), .B(Plaintext_s1[44]), .S(rst), 
        .Z(signal_1573) );
  MUX2_X1 cell_45_Ins_0_U1 ( .A(signal_794), .B(Plaintext_s0[45]), .S(rst), 
        .Z(signal_858) );
  MUX2_X1 cell_45_Ins_1_U1 ( .A(signal_1438), .B(Plaintext_s1[45]), .S(rst), 
        .Z(signal_1575) );
  MUX2_X1 cell_46_Ins_0_U1 ( .A(signal_793), .B(Plaintext_s0[46]), .S(rst), 
        .Z(signal_857) );
  MUX2_X1 cell_46_Ins_1_U1 ( .A(signal_1437), .B(Plaintext_s1[46]), .S(rst), 
        .Z(signal_1577) );
  MUX2_X1 cell_47_Ins_0_U1 ( .A(signal_792), .B(Plaintext_s0[47]), .S(rst), 
        .Z(signal_856) );
  MUX2_X1 cell_47_Ins_1_U1 ( .A(signal_1436), .B(Plaintext_s1[47]), .S(rst), 
        .Z(signal_1579) );
  MUX2_X1 cell_48_Ins_0_U1 ( .A(signal_791), .B(Plaintext_s0[48]), .S(rst), 
        .Z(signal_855) );
  MUX2_X1 cell_48_Ins_1_U1 ( .A(signal_1435), .B(Plaintext_s1[48]), .S(rst), 
        .Z(signal_1581) );
  MUX2_X1 cell_49_Ins_0_U1 ( .A(signal_790), .B(Plaintext_s0[49]), .S(rst), 
        .Z(signal_854) );
  MUX2_X1 cell_49_Ins_1_U1 ( .A(signal_1434), .B(Plaintext_s1[49]), .S(rst), 
        .Z(signal_1583) );
  MUX2_X1 cell_50_Ins_0_U1 ( .A(signal_789), .B(Plaintext_s0[50]), .S(rst), 
        .Z(signal_853) );
  MUX2_X1 cell_50_Ins_1_U1 ( .A(signal_1433), .B(Plaintext_s1[50]), .S(rst), 
        .Z(signal_1585) );
  MUX2_X1 cell_51_Ins_0_U1 ( .A(signal_788), .B(Plaintext_s0[51]), .S(rst), 
        .Z(signal_852) );
  MUX2_X1 cell_51_Ins_1_U1 ( .A(signal_1432), .B(Plaintext_s1[51]), .S(rst), 
        .Z(signal_1587) );
  MUX2_X1 cell_52_Ins_0_U1 ( .A(signal_787), .B(Plaintext_s0[52]), .S(rst), 
        .Z(signal_851) );
  MUX2_X1 cell_52_Ins_1_U1 ( .A(signal_1431), .B(Plaintext_s1[52]), .S(rst), 
        .Z(signal_1589) );
  MUX2_X1 cell_53_Ins_0_U1 ( .A(signal_786), .B(Plaintext_s0[53]), .S(rst), 
        .Z(signal_850) );
  MUX2_X1 cell_53_Ins_1_U1 ( .A(signal_1430), .B(Plaintext_s1[53]), .S(rst), 
        .Z(signal_1591) );
  MUX2_X1 cell_54_Ins_0_U1 ( .A(signal_785), .B(Plaintext_s0[54]), .S(rst), 
        .Z(signal_849) );
  MUX2_X1 cell_54_Ins_1_U1 ( .A(signal_1429), .B(Plaintext_s1[54]), .S(rst), 
        .Z(signal_1593) );
  MUX2_X1 cell_55_Ins_0_U1 ( .A(signal_784), .B(Plaintext_s0[55]), .S(rst), 
        .Z(signal_848) );
  MUX2_X1 cell_55_Ins_1_U1 ( .A(signal_1428), .B(Plaintext_s1[55]), .S(rst), 
        .Z(signal_1595) );
  MUX2_X1 cell_56_Ins_0_U1 ( .A(signal_783), .B(Plaintext_s0[56]), .S(rst), 
        .Z(signal_847) );
  MUX2_X1 cell_56_Ins_1_U1 ( .A(signal_1427), .B(Plaintext_s1[56]), .S(rst), 
        .Z(signal_1597) );
  MUX2_X1 cell_57_Ins_0_U1 ( .A(signal_782), .B(Plaintext_s0[57]), .S(rst), 
        .Z(signal_846) );
  MUX2_X1 cell_57_Ins_1_U1 ( .A(signal_1426), .B(Plaintext_s1[57]), .S(rst), 
        .Z(signal_1599) );
  MUX2_X1 cell_58_Ins_0_U1 ( .A(signal_781), .B(Plaintext_s0[58]), .S(rst), 
        .Z(signal_845) );
  MUX2_X1 cell_58_Ins_1_U1 ( .A(signal_1425), .B(Plaintext_s1[58]), .S(rst), 
        .Z(signal_1601) );
  MUX2_X1 cell_59_Ins_0_U1 ( .A(signal_780), .B(Plaintext_s0[59]), .S(rst), 
        .Z(signal_844) );
  MUX2_X1 cell_59_Ins_1_U1 ( .A(signal_1424), .B(Plaintext_s1[59]), .S(rst), 
        .Z(signal_1603) );
  MUX2_X1 cell_60_Ins_0_U1 ( .A(signal_779), .B(Plaintext_s0[60]), .S(rst), 
        .Z(signal_843) );
  MUX2_X1 cell_60_Ins_1_U1 ( .A(signal_1423), .B(Plaintext_s1[60]), .S(rst), 
        .Z(signal_1605) );
  MUX2_X1 cell_61_Ins_0_U1 ( .A(signal_778), .B(Plaintext_s0[61]), .S(rst), 
        .Z(signal_842) );
  MUX2_X1 cell_61_Ins_1_U1 ( .A(signal_1422), .B(Plaintext_s1[61]), .S(rst), 
        .Z(signal_1607) );
  MUX2_X1 cell_62_Ins_0_U1 ( .A(signal_777), .B(Plaintext_s0[62]), .S(rst), 
        .Z(signal_841) );
  MUX2_X1 cell_62_Ins_1_U1 ( .A(signal_1421), .B(Plaintext_s1[62]), .S(rst), 
        .Z(signal_1609) );
  MUX2_X1 cell_63_Ins_0_U1 ( .A(signal_776), .B(Plaintext_s0[63]), .S(rst), 
        .Z(signal_840) );
  MUX2_X1 cell_63_Ins_1_U1 ( .A(signal_1420), .B(Plaintext_s1[63]), .S(rst), 
        .Z(signal_1611) );
  XOR2_X1 cell_1000_U304 ( .A(cell_1000_n176), .B(signal_1476), .Z(signal_1428) );
  XOR2_X1 cell_1000_U303 ( .A(cell_1000_g13_1_2_), .B(signal_1475), .Z(
        signal_1427) );
  XNOR2_X1 cell_1000_U302 ( .A(cell_1000_g5_1_2_), .B(cell_1000_n175), .ZN(
        signal_1475) );
  XOR2_X1 cell_1000_U301 ( .A(1'b0), .B(cell_1000_n174), .Z(signal_1471) );
  XNOR2_X1 cell_1000_U300 ( .A(1'b0), .B(cell_1000_n173), .ZN(signal_1470) );
  XOR2_X1 cell_1000_U299 ( .A(cell_1000_n172), .B(signal_1472), .Z(signal_1424) );
  XOR2_X1 cell_1000_U298 ( .A(cell_1000_n171), .B(1'b0), .Z(signal_1469) );
  XNOR2_X1 cell_1000_U297 ( .A(1'b0), .B(cell_1000_n170), .ZN(signal_1468) );
  XNOR2_X1 cell_1000_U296 ( .A(cell_1000_n169), .B(signal_1176), .ZN(
        signal_1467) );
  XNOR2_X1 cell_1000_U295 ( .A(cell_1000_g3_1_2_), .B(cell_1000_g6_1_2_), .ZN(
        cell_1000_n169) );
  XNOR2_X1 cell_1000_U294 ( .A(cell_1000_n168), .B(cell_1000_n167), .ZN(
        signal_1466) );
  XNOR2_X1 cell_1000_U293 ( .A(cell_1000_n166), .B(cell_1000_g6_1_2_), .ZN(
        cell_1000_n167) );
  XOR2_X1 cell_1000_U292 ( .A(cell_1000_g6_1_1_), .B(signal_1179), .Z(
        cell_1000_n168) );
  XNOR2_X1 cell_1000_U291 ( .A(cell_1000_n165), .B(cell_1000_n164), .ZN(
        signal_1465) );
  XNOR2_X1 cell_1000_U290 ( .A(cell_1000_n163), .B(cell_1000_n162), .ZN(
        cell_1000_n164) );
  XNOR2_X1 cell_1000_U289 ( .A(cell_1000_g6_1_0_), .B(signal_1182), .ZN(
        cell_1000_n163) );
  XNOR2_X1 cell_1000_U288 ( .A(cell_1000_n161), .B(cell_1000_n162), .ZN(
        signal_1464) );
  XNOR2_X1 cell_1000_U287 ( .A(cell_1000_g6_1_2_), .B(cell_1000_g6_1_3_), .ZN(
        cell_1000_n162) );
  XNOR2_X1 cell_1000_U286 ( .A(signal_1185), .B(cell_1000_n160), .ZN(
        cell_1000_n161) );
  XNOR2_X1 cell_1000_U285 ( .A(cell_1000_n159), .B(signal_1188), .ZN(
        signal_1463) );
  XNOR2_X1 cell_1000_U284 ( .A(cell_1000_g4_1_2_), .B(cell_1000_g7_1_2_), .ZN(
        cell_1000_n159) );
  XNOR2_X1 cell_1000_U283 ( .A(cell_1000_n158), .B(cell_1000_n157), .ZN(
        signal_1462) );
  XNOR2_X1 cell_1000_U282 ( .A(cell_1000_n156), .B(cell_1000_g7_1_2_), .ZN(
        cell_1000_n157) );
  XOR2_X1 cell_1000_U281 ( .A(cell_1000_g7_1_1_), .B(signal_1191), .Z(
        cell_1000_n158) );
  XNOR2_X1 cell_1000_U280 ( .A(cell_1000_n155), .B(cell_1000_n154), .ZN(
        signal_1461) );
  XNOR2_X1 cell_1000_U279 ( .A(cell_1000_n153), .B(cell_1000_n152), .ZN(
        cell_1000_n154) );
  XNOR2_X1 cell_1000_U278 ( .A(cell_1000_g7_1_0_), .B(signal_1194), .ZN(
        cell_1000_n153) );
  XNOR2_X1 cell_1000_U277 ( .A(cell_1000_n151), .B(cell_1000_n152), .ZN(
        signal_1460) );
  XNOR2_X1 cell_1000_U276 ( .A(cell_1000_g7_1_2_), .B(cell_1000_g7_1_3_), .ZN(
        cell_1000_n152) );
  XNOR2_X1 cell_1000_U275 ( .A(signal_1197), .B(cell_1000_n150), .ZN(
        cell_1000_n151) );
  XNOR2_X1 cell_1000_U274 ( .A(cell_1000_n174), .B(cell_1000_n149), .ZN(
        signal_1423) );
  XOR2_X1 cell_1000_U273 ( .A(cell_1000_g8_1_2_), .B(signal_1439), .Z(
        cell_1000_n174) );
  XNOR2_X1 cell_1000_U272 ( .A(cell_1000_n148), .B(cell_1000_n147), .ZN(
        signal_1459) );
  XNOR2_X1 cell_1000_U271 ( .A(cell_1000_g5_1_2_), .B(cell_1000_n146), .ZN(
        cell_1000_n147) );
  XOR2_X1 cell_1000_U270 ( .A(1'b0), .B(signal_1200), .Z(cell_1000_n148) );
  XOR2_X1 cell_1000_U269 ( .A(cell_1000_n145), .B(cell_1000_n144), .Z(
        signal_1458) );
  XNOR2_X1 cell_1000_U268 ( .A(cell_1000_n143), .B(cell_1000_n142), .ZN(
        cell_1000_n144) );
  XNOR2_X1 cell_1000_U267 ( .A(cell_1000_n146), .B(cell_1000_g14_1_1_), .ZN(
        cell_1000_n142) );
  XOR2_X1 cell_1000_U266 ( .A(1'b0), .B(cell_1000_g14_1_2_), .Z(cell_1000_n146) );
  XOR2_X1 cell_1000_U265 ( .A(1'b0), .B(signal_1203), .Z(cell_1000_n143) );
  XNOR2_X1 cell_1000_U264 ( .A(cell_1000_n141), .B(cell_1000_n140), .ZN(
        signal_1457) );
  XNOR2_X1 cell_1000_U263 ( .A(cell_1000_n139), .B(cell_1000_n138), .ZN(
        cell_1000_n140) );
  XNOR2_X1 cell_1000_U262 ( .A(cell_1000_g14_1_0_), .B(signal_1206), .ZN(
        cell_1000_n139) );
  XNOR2_X1 cell_1000_U261 ( .A(cell_1000_n137), .B(cell_1000_n138), .ZN(
        signal_1456) );
  XNOR2_X1 cell_1000_U260 ( .A(cell_1000_g14_1_2_), .B(cell_1000_g14_1_3_), 
        .ZN(cell_1000_n138) );
  XNOR2_X1 cell_1000_U259 ( .A(signal_1209), .B(cell_1000_n136), .ZN(
        cell_1000_n137) );
  XNOR2_X1 cell_1000_U258 ( .A(cell_1000_n135), .B(signal_1164), .ZN(
        signal_1455) );
  XNOR2_X1 cell_1000_U257 ( .A(cell_1000_g8_1_2_), .B(cell_1000_g9_1_2_), .ZN(
        cell_1000_n135) );
  XNOR2_X1 cell_1000_U256 ( .A(cell_1000_n134), .B(cell_1000_n133), .ZN(
        signal_1454) );
  XNOR2_X1 cell_1000_U255 ( .A(cell_1000_n132), .B(cell_1000_g9_1_2_), .ZN(
        cell_1000_n133) );
  XOR2_X1 cell_1000_U254 ( .A(cell_1000_g9_1_1_), .B(signal_1167), .Z(
        cell_1000_n134) );
  XNOR2_X1 cell_1000_U253 ( .A(cell_1000_n131), .B(cell_1000_n130), .ZN(
        signal_1453) );
  XNOR2_X1 cell_1000_U252 ( .A(cell_1000_n129), .B(cell_1000_n128), .ZN(
        cell_1000_n130) );
  XNOR2_X1 cell_1000_U251 ( .A(cell_1000_g9_1_0_), .B(signal_1170), .ZN(
        cell_1000_n131) );
  XNOR2_X1 cell_1000_U250 ( .A(cell_1000_n127), .B(signal_1173), .ZN(
        signal_1452) );
  XNOR2_X1 cell_1000_U249 ( .A(cell_1000_n126), .B(cell_1000_n128), .ZN(
        cell_1000_n127) );
  XOR2_X1 cell_1000_U248 ( .A(cell_1000_g9_1_2_), .B(cell_1000_g9_1_3_), .Z(
        cell_1000_n128) );
  XNOR2_X1 cell_1000_U247 ( .A(1'b0), .B(cell_1000_n125), .ZN(signal_1451) );
  XNOR2_X1 cell_1000_U246 ( .A(1'b0), .B(cell_1000_n124), .ZN(signal_1450) );
  XNOR2_X1 cell_1000_U245 ( .A(cell_1000_n123), .B(cell_1000_n173), .ZN(
        signal_1422) );
  XNOR2_X1 cell_1000_U244 ( .A(signal_1438), .B(cell_1000_n132), .ZN(
        cell_1000_n173) );
  XOR2_X1 cell_1000_U243 ( .A(cell_1000_g8_1_2_), .B(cell_1000_g8_1_1_), .Z(
        cell_1000_n132) );
  XNOR2_X1 cell_1000_U242 ( .A(cell_1000_g15_1[1]), .B(cell_1000_n149), .ZN(
        cell_1000_n123) );
  XNOR2_X1 cell_1000_U241 ( .A(1'b0), .B(cell_1000_n122), .ZN(signal_1449) );
  XNOR2_X1 cell_1000_U240 ( .A(1'b0), .B(cell_1000_n121), .ZN(signal_1447) );
  XNOR2_X1 cell_1000_U239 ( .A(1'b0), .B(cell_1000_n120), .ZN(signal_1446) );
  XNOR2_X1 cell_1000_U238 ( .A(1'b0), .B(cell_1000_n119), .ZN(signal_1445) );
  XNOR2_X1 cell_1000_U237 ( .A(1'b0), .B(cell_1000_n175), .ZN(signal_1443) );
  XNOR2_X1 cell_1000_U236 ( .A(cell_1000_g2_1_2_), .B(signal_1236), .ZN(
        cell_1000_n175) );
  XNOR2_X1 cell_1000_U235 ( .A(1'b0), .B(cell_1000_n118), .ZN(signal_1442) );
  XNOR2_X1 cell_1000_U234 ( .A(1'b0), .B(cell_1000_n117), .ZN(signal_1441) );
  XNOR2_X1 cell_1000_U233 ( .A(cell_1000_n116), .B(cell_1000_n115), .ZN(
        signal_1421) );
  XNOR2_X1 cell_1000_U232 ( .A(cell_1000_n171), .B(cell_1000_g15_1[0]), .ZN(
        cell_1000_n116) );
  XNOR2_X1 cell_1000_U231 ( .A(signal_1437), .B(cell_1000_n129), .ZN(
        cell_1000_n171) );
  XNOR2_X1 cell_1000_U230 ( .A(cell_1000_g8_1_0_), .B(cell_1000_n126), .ZN(
        cell_1000_n129) );
  XNOR2_X1 cell_1000_U229 ( .A(cell_1000_n114), .B(signal_1248), .ZN(
        signal_1439) );
  XNOR2_X1 cell_1000_U228 ( .A(cell_1000_g10_1_2_), .B(1'b0), .ZN(
        cell_1000_n114) );
  XNOR2_X1 cell_1000_U227 ( .A(cell_1000_n113), .B(cell_1000_n112), .ZN(
        signal_1438) );
  XNOR2_X1 cell_1000_U226 ( .A(cell_1000_g10_1_2_), .B(1'b0), .ZN(
        cell_1000_n112) );
  XOR2_X1 cell_1000_U225 ( .A(cell_1000_g10_1_1_), .B(signal_1251), .Z(
        cell_1000_n113) );
  XNOR2_X1 cell_1000_U224 ( .A(cell_1000_n111), .B(cell_1000_n110), .ZN(
        signal_1437) );
  XNOR2_X1 cell_1000_U223 ( .A(cell_1000_n109), .B(signal_1254), .ZN(
        cell_1000_n110) );
  XOR2_X1 cell_1000_U222 ( .A(1'b0), .B(cell_1000_g10_1_0_), .Z(cell_1000_n111) );
  XOR2_X1 cell_1000_U221 ( .A(cell_1000_g11_1_2_), .B(signal_1483), .Z(
        signal_1435) );
  XNOR2_X1 cell_1000_U220 ( .A(cell_1000_g3_1_2_), .B(cell_1000_n125), .ZN(
        signal_1483) );
  XNOR2_X1 cell_1000_U219 ( .A(cell_1000_g0_1_2_), .B(signal_1212), .ZN(
        cell_1000_n125) );
  XOR2_X1 cell_1000_U218 ( .A(cell_1000_n108), .B(signal_1480), .Z(signal_1432) );
  XNOR2_X1 cell_1000_U217 ( .A(cell_1000_n107), .B(cell_1000_n160), .ZN(
        signal_1480) );
  XOR2_X1 cell_1000_U216 ( .A(cell_1000_g12_1_2_), .B(signal_1479), .Z(
        signal_1431) );
  XNOR2_X1 cell_1000_U215 ( .A(cell_1000_g4_1_2_), .B(cell_1000_n121), .ZN(
        signal_1479) );
  XNOR2_X1 cell_1000_U214 ( .A(cell_1000_g1_1_2_), .B(signal_1224), .ZN(
        cell_1000_n121) );
  XNOR2_X1 cell_1000_U213 ( .A(cell_1000_n115), .B(cell_1000_n170), .ZN(
        signal_1420) );
  XNOR2_X1 cell_1000_U212 ( .A(cell_1000_n126), .B(signal_1436), .ZN(
        cell_1000_n170) );
  XOR2_X1 cell_1000_U211 ( .A(cell_1000_g8_1_2_), .B(cell_1000_g8_1_3_), .Z(
        cell_1000_n126) );
  XNOR2_X1 cell_1000_U210 ( .A(cell_1000_g15_1[3]), .B(cell_1000_n149), .ZN(
        cell_1000_n115) );
  XNOR2_X1 cell_1000_U209 ( .A(1'b0), .B(cell_1000_g15_1[2]), .ZN(
        cell_1000_n149) );
  XNOR2_X1 cell_1000_U208 ( .A(cell_1000_g12_0_0_), .B(cell_1000_n106), .ZN(
        signal_785) );
  XOR2_X1 cell_1000_U207 ( .A(cell_1000_n105), .B(signal_833), .Z(
        cell_1000_n106) );
  XNOR2_X1 cell_1000_U206 ( .A(cell_1000_n105), .B(signal_832), .ZN(signal_784) );
  XOR2_X1 cell_1000_U205 ( .A(cell_1000_g12_0_2_), .B(cell_1000_g12_0_3_), .Z(
        cell_1000_n105) );
  XOR2_X1 cell_1000_U204 ( .A(cell_1000_g13_0_2_), .B(signal_831), .Z(
        signal_783) );
  XNOR2_X1 cell_1000_U203 ( .A(cell_1000_g13_0_0_), .B(cell_1000_n104), .ZN(
        signal_781) );
  XOR2_X1 cell_1000_U202 ( .A(cell_1000_n103), .B(signal_829), .Z(
        cell_1000_n104) );
  XNOR2_X1 cell_1000_U201 ( .A(cell_1000_n102), .B(cell_1000_n101), .ZN(
        signal_833) );
  XNOR2_X1 cell_1000_U200 ( .A(cell_1000_n100), .B(cell_1000_n99), .ZN(
        signal_832) );
  XNOR2_X1 cell_1000_U199 ( .A(cell_1000_g5_0_2_), .B(cell_1000_n98), .ZN(
        signal_831) );
  XNOR2_X1 cell_1000_U198 ( .A(cell_1000_n97), .B(cell_1000_n96), .ZN(
        signal_829) );
  XNOR2_X1 cell_1000_U197 ( .A(1'b0), .B(cell_1000_n95), .ZN(signal_827) );
  XOR2_X1 cell_1000_U196 ( .A(1'b0), .B(cell_1000_n94), .Z(signal_826) );
  XNOR2_X1 cell_1000_U195 ( .A(cell_1000_n103), .B(signal_828), .ZN(signal_780) );
  XOR2_X1 cell_1000_U194 ( .A(cell_1000_g13_0_2_), .B(cell_1000_g13_0_3_), .Z(
        cell_1000_n103) );
  XNOR2_X1 cell_1000_U193 ( .A(cell_1000_n93), .B(cell_1000_n92), .ZN(
        signal_828) );
  XOR2_X1 cell_1000_U192 ( .A(cell_1000_n91), .B(1'b0), .Z(signal_825) );
  XNOR2_X1 cell_1000_U191 ( .A(1'b0), .B(cell_1000_n90), .ZN(signal_824) );
  XNOR2_X1 cell_1000_U190 ( .A(cell_1000_n89), .B(signal_1159), .ZN(signal_823) );
  XNOR2_X1 cell_1000_U189 ( .A(cell_1000_g3_0_2_), .B(cell_1000_g6_0_2_), .ZN(
        cell_1000_n89) );
  XNOR2_X1 cell_1000_U188 ( .A(cell_1000_n88), .B(cell_1000_n87), .ZN(
        signal_822) );
  XNOR2_X1 cell_1000_U187 ( .A(cell_1000_n86), .B(cell_1000_g6_0_2_), .ZN(
        cell_1000_n87) );
  XOR2_X1 cell_1000_U186 ( .A(cell_1000_g6_0_1_), .B(signal_1158), .Z(
        cell_1000_n88) );
  XNOR2_X1 cell_1000_U185 ( .A(cell_1000_n85), .B(cell_1000_n84), .ZN(
        signal_821) );
  XNOR2_X1 cell_1000_U184 ( .A(cell_1000_n83), .B(cell_1000_n82), .ZN(
        cell_1000_n84) );
  XOR2_X1 cell_1000_U183 ( .A(signal_1157), .B(cell_1000_g6_0_0_), .Z(
        cell_1000_n85) );
  XNOR2_X1 cell_1000_U182 ( .A(cell_1000_n81), .B(signal_1156), .ZN(signal_820) );
  XNOR2_X1 cell_1000_U181 ( .A(cell_1000_n80), .B(cell_1000_n82), .ZN(
        cell_1000_n81) );
  XOR2_X1 cell_1000_U180 ( .A(cell_1000_g6_0_2_), .B(cell_1000_g6_0_3_), .Z(
        cell_1000_n82) );
  XNOR2_X1 cell_1000_U179 ( .A(cell_1000_n79), .B(signal_1155), .ZN(signal_819) );
  XNOR2_X1 cell_1000_U178 ( .A(cell_1000_g4_0_2_), .B(cell_1000_g7_0_2_), .ZN(
        cell_1000_n79) );
  XNOR2_X1 cell_1000_U177 ( .A(cell_1000_n78), .B(cell_1000_n77), .ZN(
        signal_818) );
  XNOR2_X1 cell_1000_U176 ( .A(cell_1000_n76), .B(signal_1154), .ZN(
        cell_1000_n77) );
  XNOR2_X1 cell_1000_U175 ( .A(cell_1000_g7_0_2_), .B(cell_1000_g7_0_1_), .ZN(
        cell_1000_n76) );
  XNOR2_X1 cell_1000_U174 ( .A(cell_1000_n75), .B(cell_1000_n74), .ZN(
        signal_817) );
  XNOR2_X1 cell_1000_U173 ( .A(cell_1000_n102), .B(cell_1000_n73), .ZN(
        cell_1000_n74) );
  XOR2_X1 cell_1000_U172 ( .A(cell_1000_n100), .B(cell_1000_g4_0_0_), .Z(
        cell_1000_n102) );
  XOR2_X1 cell_1000_U171 ( .A(signal_1153), .B(cell_1000_g7_0_0_), .Z(
        cell_1000_n75) );
  XNOR2_X1 cell_1000_U170 ( .A(cell_1000_n72), .B(signal_1152), .ZN(signal_816) );
  XNOR2_X1 cell_1000_U169 ( .A(cell_1000_n100), .B(cell_1000_n73), .ZN(
        cell_1000_n72) );
  XOR2_X1 cell_1000_U168 ( .A(cell_1000_g7_0_2_), .B(cell_1000_g7_0_3_), .Z(
        cell_1000_n73) );
  XOR2_X1 cell_1000_U167 ( .A(cell_1000_g4_0_2_), .B(cell_1000_g4_0_3_), .Z(
        cell_1000_n100) );
  XNOR2_X1 cell_1000_U166 ( .A(cell_1000_n71), .B(cell_1000_n95), .ZN(
        signal_779) );
  XNOR2_X1 cell_1000_U165 ( .A(cell_1000_g8_0_2_), .B(signal_795), .ZN(
        cell_1000_n95) );
  XNOR2_X1 cell_1000_U164 ( .A(cell_1000_n70), .B(cell_1000_n69), .ZN(
        signal_815) );
  XNOR2_X1 cell_1000_U163 ( .A(cell_1000_g5_0_2_), .B(cell_1000_n68), .ZN(
        cell_1000_n69) );
  XOR2_X1 cell_1000_U162 ( .A(signal_940), .B(signal_1151), .Z(cell_1000_n70)
         );
  XOR2_X1 cell_1000_U161 ( .A(cell_1000_n67), .B(cell_1000_n66), .Z(signal_814) );
  XNOR2_X1 cell_1000_U160 ( .A(cell_1000_n65), .B(cell_1000_n64), .ZN(
        cell_1000_n66) );
  XNOR2_X1 cell_1000_U159 ( .A(cell_1000_n68), .B(cell_1000_g14_0_1_), .ZN(
        cell_1000_n64) );
  XOR2_X1 cell_1000_U158 ( .A(1'b0), .B(cell_1000_g14_0_2_), .Z(cell_1000_n68)
         );
  XOR2_X1 cell_1000_U157 ( .A(signal_939), .B(signal_1150), .Z(cell_1000_n65)
         );
  XNOR2_X1 cell_1000_U156 ( .A(cell_1000_n63), .B(cell_1000_n62), .ZN(
        signal_813) );
  XNOR2_X1 cell_1000_U155 ( .A(cell_1000_n97), .B(cell_1000_n61), .ZN(
        cell_1000_n62) );
  XOR2_X1 cell_1000_U154 ( .A(cell_1000_n93), .B(cell_1000_g5_0_0_), .Z(
        cell_1000_n97) );
  XOR2_X1 cell_1000_U153 ( .A(signal_1149), .B(cell_1000_g14_0_0_), .Z(
        cell_1000_n63) );
  XNOR2_X1 cell_1000_U152 ( .A(cell_1000_n60), .B(signal_1148), .ZN(signal_812) );
  XNOR2_X1 cell_1000_U151 ( .A(cell_1000_n93), .B(cell_1000_n61), .ZN(
        cell_1000_n60) );
  XOR2_X1 cell_1000_U150 ( .A(cell_1000_g14_0_2_), .B(cell_1000_g14_0_3_), .Z(
        cell_1000_n61) );
  XOR2_X1 cell_1000_U149 ( .A(cell_1000_g5_0_2_), .B(cell_1000_g5_0_3_), .Z(
        cell_1000_n93) );
  XNOR2_X1 cell_1000_U148 ( .A(cell_1000_n59), .B(signal_1163), .ZN(signal_811) );
  XNOR2_X1 cell_1000_U147 ( .A(cell_1000_g8_0_2_), .B(cell_1000_g9_0_2_), .ZN(
        cell_1000_n59) );
  XNOR2_X1 cell_1000_U146 ( .A(cell_1000_n58), .B(cell_1000_n57), .ZN(
        signal_810) );
  XNOR2_X1 cell_1000_U145 ( .A(cell_1000_n56), .B(cell_1000_g9_0_2_), .ZN(
        cell_1000_n57) );
  XNOR2_X1 cell_1000_U144 ( .A(signal_1162), .B(cell_1000_g9_0_1_), .ZN(
        cell_1000_n58) );
  XNOR2_X1 cell_1000_U143 ( .A(cell_1000_n55), .B(cell_1000_n54), .ZN(
        signal_809) );
  XNOR2_X1 cell_1000_U142 ( .A(cell_1000_n53), .B(cell_1000_n52), .ZN(
        cell_1000_n54) );
  XNOR2_X1 cell_1000_U141 ( .A(signal_1161), .B(cell_1000_g9_0_0_), .ZN(
        cell_1000_n53) );
  XNOR2_X1 cell_1000_U140 ( .A(cell_1000_n51), .B(cell_1000_n52), .ZN(
        signal_808) );
  XNOR2_X1 cell_1000_U139 ( .A(cell_1000_g9_0_2_), .B(cell_1000_g9_0_3_), .ZN(
        cell_1000_n52) );
  XNOR2_X1 cell_1000_U138 ( .A(signal_1160), .B(cell_1000_n50), .ZN(
        cell_1000_n51) );
  XNOR2_X1 cell_1000_U137 ( .A(1'b0), .B(cell_1000_n49), .ZN(signal_807) );
  XNOR2_X1 cell_1000_U136 ( .A(1'b0), .B(cell_1000_n48), .ZN(signal_806) );
  XNOR2_X1 cell_1000_U135 ( .A(cell_1000_n47), .B(cell_1000_g15_0[1]), .ZN(
        signal_778) );
  XNOR2_X1 cell_1000_U134 ( .A(cell_1000_n71), .B(cell_1000_n94), .ZN(
        cell_1000_n47) );
  XNOR2_X1 cell_1000_U133 ( .A(signal_794), .B(cell_1000_n56), .ZN(
        cell_1000_n94) );
  XNOR2_X1 cell_1000_U132 ( .A(cell_1000_g8_0_2_), .B(cell_1000_g8_0_1_), .ZN(
        cell_1000_n56) );
  XOR2_X1 cell_1000_U131 ( .A(1'b0), .B(cell_1000_n46), .Z(signal_805) );
  XOR2_X1 cell_1000_U130 ( .A(1'b0), .B(cell_1000_n45), .Z(signal_804) );
  XOR2_X1 cell_1000_U129 ( .A(1'b0), .B(cell_1000_n44), .Z(signal_802) );
  XOR2_X1 cell_1000_U128 ( .A(1'b0), .B(cell_1000_n101), .Z(signal_801) );
  XNOR2_X1 cell_1000_U127 ( .A(cell_1000_g1_0_0_), .B(cell_1000_n43), .ZN(
        cell_1000_n101) );
  XOR2_X1 cell_1000_U126 ( .A(cell_1000_n42), .B(signal_1141), .Z(
        cell_1000_n43) );
  XOR2_X1 cell_1000_U125 ( .A(1'b0), .B(cell_1000_n99), .Z(signal_800) );
  XNOR2_X1 cell_1000_U124 ( .A(cell_1000_n42), .B(signal_1140), .ZN(
        cell_1000_n99) );
  XOR2_X1 cell_1000_U123 ( .A(cell_1000_g1_0_2_), .B(cell_1000_g1_0_3_), .Z(
        cell_1000_n42) );
  XNOR2_X1 cell_1000_U122 ( .A(1'b0), .B(cell_1000_n98), .ZN(signal_799) );
  XNOR2_X1 cell_1000_U121 ( .A(cell_1000_g2_0_2_), .B(signal_1139), .ZN(
        cell_1000_n98) );
  XNOR2_X1 cell_1000_U120 ( .A(1'b0), .B(cell_1000_n41), .ZN(signal_798) );
  XOR2_X1 cell_1000_U119 ( .A(1'b0), .B(cell_1000_n96), .Z(signal_797) );
  XNOR2_X1 cell_1000_U118 ( .A(cell_1000_g2_0_0_), .B(cell_1000_n40), .ZN(
        cell_1000_n96) );
  XOR2_X1 cell_1000_U117 ( .A(cell_1000_n39), .B(signal_1137), .Z(
        cell_1000_n40) );
  XOR2_X1 cell_1000_U116 ( .A(1'b0), .B(cell_1000_n92), .Z(signal_796) );
  XNOR2_X1 cell_1000_U115 ( .A(cell_1000_n39), .B(signal_1136), .ZN(
        cell_1000_n92) );
  XOR2_X1 cell_1000_U114 ( .A(cell_1000_g2_0_2_), .B(cell_1000_g2_0_3_), .Z(
        cell_1000_n39) );
  XNOR2_X1 cell_1000_U113 ( .A(cell_1000_n38), .B(cell_1000_n37), .ZN(
        signal_777) );
  XNOR2_X1 cell_1000_U112 ( .A(cell_1000_n91), .B(cell_1000_g15_0[0]), .ZN(
        cell_1000_n38) );
  XNOR2_X1 cell_1000_U111 ( .A(cell_1000_n55), .B(signal_793), .ZN(
        cell_1000_n91) );
  XNOR2_X1 cell_1000_U110 ( .A(cell_1000_g8_0_0_), .B(cell_1000_n50), .ZN(
        cell_1000_n55) );
  XNOR2_X1 cell_1000_U109 ( .A(cell_1000_n36), .B(signal_1135), .ZN(signal_795) );
  XNOR2_X1 cell_1000_U108 ( .A(cell_1000_g10_0_2_), .B(signal_1028), .ZN(
        cell_1000_n36) );
  XNOR2_X1 cell_1000_U107 ( .A(cell_1000_n35), .B(cell_1000_n34), .ZN(
        signal_794) );
  XNOR2_X1 cell_1000_U106 ( .A(cell_1000_g10_0_2_), .B(signal_943), .ZN(
        cell_1000_n34) );
  XOR2_X1 cell_1000_U105 ( .A(cell_1000_g10_0_1_), .B(signal_1134), .Z(
        cell_1000_n35) );
  XNOR2_X1 cell_1000_U104 ( .A(cell_1000_n33), .B(cell_1000_n32), .ZN(
        signal_793) );
  XNOR2_X1 cell_1000_U103 ( .A(cell_1000_n31), .B(signal_1133), .ZN(
        cell_1000_n32) );
  XNOR2_X1 cell_1000_U102 ( .A(cell_1000_g10_0_0_), .B(signal_1026), .ZN(
        cell_1000_n31) );
  XOR2_X1 cell_1000_U101 ( .A(cell_1000_g11_0_2_), .B(signal_839), .Z(
        signal_791) );
  XNOR2_X1 cell_1000_U100 ( .A(cell_1000_g3_0_2_), .B(cell_1000_n49), .ZN(
        signal_839) );
  XNOR2_X1 cell_1000_U99 ( .A(cell_1000_g0_0_2_), .B(signal_1147), .ZN(
        cell_1000_n49) );
  XNOR2_X1 cell_1000_U98 ( .A(cell_1000_g11_0_0_), .B(cell_1000_n30), .ZN(
        signal_789) );
  XOR2_X1 cell_1000_U97 ( .A(cell_1000_n29), .B(signal_837), .Z(cell_1000_n30)
         );
  XNOR2_X1 cell_1000_U96 ( .A(cell_1000_n83), .B(cell_1000_n46), .ZN(
        signal_837) );
  XNOR2_X1 cell_1000_U95 ( .A(cell_1000_g0_0_0_), .B(cell_1000_n28), .ZN(
        cell_1000_n46) );
  XOR2_X1 cell_1000_U94 ( .A(cell_1000_n27), .B(signal_1145), .Z(cell_1000_n28) );
  XOR2_X1 cell_1000_U93 ( .A(cell_1000_n80), .B(cell_1000_g3_0_0_), .Z(
        cell_1000_n83) );
  XNOR2_X1 cell_1000_U92 ( .A(cell_1000_n29), .B(signal_836), .ZN(signal_788)
         );
  XOR2_X1 cell_1000_U91 ( .A(cell_1000_g11_0_2_), .B(cell_1000_g11_0_3_), .Z(
        cell_1000_n29) );
  XNOR2_X1 cell_1000_U90 ( .A(cell_1000_n80), .B(cell_1000_n45), .ZN(
        signal_836) );
  XNOR2_X1 cell_1000_U89 ( .A(cell_1000_n27), .B(signal_1144), .ZN(
        cell_1000_n45) );
  XOR2_X1 cell_1000_U88 ( .A(cell_1000_g0_0_2_), .B(cell_1000_g0_0_3_), .Z(
        cell_1000_n27) );
  XOR2_X1 cell_1000_U87 ( .A(cell_1000_g3_0_2_), .B(cell_1000_g3_0_3_), .Z(
        cell_1000_n80) );
  XOR2_X1 cell_1000_U86 ( .A(cell_1000_g12_0_2_), .B(signal_835), .Z(
        signal_787) );
  XNOR2_X1 cell_1000_U85 ( .A(cell_1000_n26), .B(signal_834), .ZN(signal_786)
         );
  XNOR2_X1 cell_1000_U84 ( .A(cell_1000_g12_0_2_), .B(cell_1000_g12_0_1_), 
        .ZN(cell_1000_n26) );
  XNOR2_X1 cell_1000_U83 ( .A(cell_1000_n78), .B(cell_1000_n44), .ZN(
        signal_834) );
  XNOR2_X1 cell_1000_U82 ( .A(cell_1000_n25), .B(cell_1000_g1_0_1_), .ZN(
        cell_1000_n44) );
  XNOR2_X1 cell_1000_U81 ( .A(cell_1000_g1_0_2_), .B(signal_1142), .ZN(
        cell_1000_n25) );
  XOR2_X1 cell_1000_U80 ( .A(cell_1000_g4_0_2_), .B(cell_1000_g4_0_1_), .Z(
        cell_1000_n78) );
  XNOR2_X1 cell_1000_U79 ( .A(cell_1000_n37), .B(cell_1000_n90), .ZN(
        signal_776) );
  XNOR2_X1 cell_1000_U78 ( .A(cell_1000_n50), .B(signal_792), .ZN(
        cell_1000_n90) );
  XNOR2_X1 cell_1000_U77 ( .A(signal_1132), .B(cell_1000_n24), .ZN(signal_792)
         );
  XOR2_X1 cell_1000_U76 ( .A(cell_1000_n33), .B(signal_1025), .Z(cell_1000_n24) );
  XOR2_X1 cell_1000_U75 ( .A(cell_1000_g10_0_2_), .B(cell_1000_g10_0_3_), .Z(
        cell_1000_n33) );
  XNOR2_X1 cell_1000_U74 ( .A(cell_1000_g8_0_2_), .B(cell_1000_g8_0_3_), .ZN(
        cell_1000_n50) );
  XNOR2_X1 cell_1000_U73 ( .A(cell_1000_n71), .B(cell_1000_g15_0[3]), .ZN(
        cell_1000_n37) );
  XOR2_X1 cell_1000_U72 ( .A(1'b0), .B(cell_1000_g15_0[2]), .Z(cell_1000_n71)
         );
  XNOR2_X1 cell_1000_U71 ( .A(cell_1000_n23), .B(cell_1000_g11_1_0_), .ZN(
        signal_1433) );
  XNOR2_X1 cell_1000_U70 ( .A(cell_1000_n108), .B(signal_1481), .ZN(
        cell_1000_n23) );
  XOR2_X1 cell_1000_U69 ( .A(cell_1000_g11_1_2_), .B(cell_1000_g11_1_3_), .Z(
        cell_1000_n108) );
  XNOR2_X1 cell_1000_U68 ( .A(cell_1000_n165), .B(cell_1000_n122), .ZN(
        signal_1481) );
  XNOR2_X1 cell_1000_U67 ( .A(cell_1000_n22), .B(cell_1000_n21), .ZN(
        cell_1000_n122) );
  XNOR2_X1 cell_1000_U66 ( .A(signal_1218), .B(cell_1000_g0_1_0_), .ZN(
        cell_1000_n22) );
  XNOR2_X1 cell_1000_U65 ( .A(cell_1000_g3_1_0_), .B(cell_1000_n160), .ZN(
        cell_1000_n165) );
  XNOR2_X1 cell_1000_U64 ( .A(cell_1000_g3_1_2_), .B(cell_1000_g3_1_3_), .ZN(
        cell_1000_n160) );
  XNOR2_X1 cell_1000_U63 ( .A(cell_1000_n20), .B(cell_1000_g11_1_1_), .ZN(
        signal_1434) );
  XNOR2_X1 cell_1000_U62 ( .A(cell_1000_g11_1_2_), .B(signal_1482), .ZN(
        cell_1000_n20) );
  XNOR2_X1 cell_1000_U61 ( .A(cell_1000_n166), .B(cell_1000_n124), .ZN(
        signal_1482) );
  XNOR2_X1 cell_1000_U60 ( .A(cell_1000_g0_1_1_), .B(cell_1000_n19), .ZN(
        cell_1000_n124) );
  XOR2_X1 cell_1000_U59 ( .A(cell_1000_g0_1_2_), .B(signal_1215), .Z(
        cell_1000_n19) );
  XOR2_X1 cell_1000_U58 ( .A(cell_1000_g3_1_2_), .B(cell_1000_g3_1_1_), .Z(
        cell_1000_n166) );
  XOR2_X1 cell_1000_U57 ( .A(1'b0), .B(cell_1000_n107), .Z(signal_1448) );
  XNOR2_X1 cell_1000_U56 ( .A(signal_1221), .B(cell_1000_n21), .ZN(
        cell_1000_n107) );
  XNOR2_X1 cell_1000_U55 ( .A(cell_1000_g0_1_2_), .B(cell_1000_g0_1_3_), .ZN(
        cell_1000_n21) );
  XNOR2_X1 cell_1000_U54 ( .A(cell_1000_n18), .B(cell_1000_g11_0_1_), .ZN(
        signal_790) );
  XNOR2_X1 cell_1000_U53 ( .A(cell_1000_g11_0_2_), .B(signal_838), .ZN(
        cell_1000_n18) );
  XNOR2_X1 cell_1000_U52 ( .A(cell_1000_n86), .B(cell_1000_n48), .ZN(
        signal_838) );
  XNOR2_X1 cell_1000_U51 ( .A(cell_1000_g0_0_1_), .B(cell_1000_n17), .ZN(
        cell_1000_n48) );
  XOR2_X1 cell_1000_U50 ( .A(cell_1000_g0_0_2_), .B(signal_1146), .Z(
        cell_1000_n17) );
  XOR2_X1 cell_1000_U49 ( .A(cell_1000_g3_0_2_), .B(cell_1000_g3_0_1_), .Z(
        cell_1000_n86) );
  XNOR2_X1 cell_1000_U48 ( .A(cell_1000_n16), .B(cell_1000_g12_1_0_), .ZN(
        signal_1429) );
  XNOR2_X1 cell_1000_U47 ( .A(cell_1000_n176), .B(signal_1477), .ZN(
        cell_1000_n16) );
  XOR2_X1 cell_1000_U46 ( .A(cell_1000_g12_1_2_), .B(cell_1000_g12_1_3_), .Z(
        cell_1000_n176) );
  XNOR2_X1 cell_1000_U45 ( .A(cell_1000_n155), .B(cell_1000_n119), .ZN(
        signal_1477) );
  XNOR2_X1 cell_1000_U44 ( .A(cell_1000_n15), .B(cell_1000_n14), .ZN(
        cell_1000_n119) );
  XNOR2_X1 cell_1000_U43 ( .A(signal_1230), .B(cell_1000_g1_1_0_), .ZN(
        cell_1000_n15) );
  XNOR2_X1 cell_1000_U42 ( .A(cell_1000_g4_1_0_), .B(cell_1000_n150), .ZN(
        cell_1000_n155) );
  XNOR2_X1 cell_1000_U41 ( .A(cell_1000_n13), .B(cell_1000_g12_1_1_), .ZN(
        signal_1430) );
  XNOR2_X1 cell_1000_U40 ( .A(cell_1000_g12_1_2_), .B(signal_1478), .ZN(
        cell_1000_n13) );
  XNOR2_X1 cell_1000_U39 ( .A(cell_1000_n156), .B(cell_1000_n120), .ZN(
        signal_1478) );
  XNOR2_X1 cell_1000_U38 ( .A(cell_1000_g1_1_1_), .B(cell_1000_n12), .ZN(
        cell_1000_n120) );
  XOR2_X1 cell_1000_U37 ( .A(cell_1000_g1_1_2_), .B(signal_1227), .Z(
        cell_1000_n12) );
  XOR2_X1 cell_1000_U36 ( .A(cell_1000_g4_1_2_), .B(cell_1000_g4_1_1_), .Z(
        cell_1000_n156) );
  XOR2_X1 cell_1000_U35 ( .A(1'b0), .B(cell_1000_n11), .Z(signal_1444) );
  XNOR2_X1 cell_1000_U34 ( .A(1'b0), .B(cell_1000_n10), .ZN(signal_803) );
  XNOR2_X1 cell_1000_U33 ( .A(cell_1000_n9), .B(cell_1000_g13_1_0_), .ZN(
        signal_1425) );
  XNOR2_X1 cell_1000_U32 ( .A(cell_1000_n172), .B(signal_1473), .ZN(
        cell_1000_n9) );
  XOR2_X1 cell_1000_U31 ( .A(cell_1000_g13_1_2_), .B(cell_1000_g13_1_3_), .Z(
        cell_1000_n172) );
  XNOR2_X1 cell_1000_U30 ( .A(cell_1000_n141), .B(cell_1000_n117), .ZN(
        signal_1473) );
  XNOR2_X1 cell_1000_U29 ( .A(cell_1000_n8), .B(cell_1000_n7), .ZN(
        cell_1000_n117) );
  XNOR2_X1 cell_1000_U28 ( .A(signal_1242), .B(cell_1000_g2_1_0_), .ZN(
        cell_1000_n8) );
  XNOR2_X1 cell_1000_U27 ( .A(cell_1000_g5_1_0_), .B(cell_1000_n136), .ZN(
        cell_1000_n141) );
  XNOR2_X1 cell_1000_U26 ( .A(cell_1000_n6), .B(cell_1000_g13_1_1_), .ZN(
        signal_1426) );
  XNOR2_X1 cell_1000_U25 ( .A(cell_1000_g13_1_2_), .B(signal_1474), .ZN(
        cell_1000_n6) );
  XNOR2_X1 cell_1000_U24 ( .A(cell_1000_n145), .B(cell_1000_n118), .ZN(
        signal_1474) );
  XNOR2_X1 cell_1000_U23 ( .A(signal_1239), .B(cell_1000_n5), .ZN(
        cell_1000_n118) );
  XOR2_X1 cell_1000_U22 ( .A(cell_1000_g2_1_2_), .B(cell_1000_g2_1_1_), .Z(
        cell_1000_n5) );
  XOR2_X1 cell_1000_U21 ( .A(cell_1000_g5_1_2_), .B(cell_1000_g5_1_1_), .Z(
        cell_1000_n145) );
  XOR2_X1 cell_1000_U20 ( .A(1'b0), .B(cell_1000_n4), .Z(signal_1440) );
  XNOR2_X1 cell_1000_U19 ( .A(cell_1000_n3), .B(cell_1000_g13_0_1_), .ZN(
        signal_782) );
  XNOR2_X1 cell_1000_U18 ( .A(cell_1000_g13_0_2_), .B(signal_830), .ZN(
        cell_1000_n3) );
  XNOR2_X1 cell_1000_U17 ( .A(cell_1000_n67), .B(cell_1000_n41), .ZN(
        signal_830) );
  XNOR2_X1 cell_1000_U16 ( .A(signal_1138), .B(cell_1000_n2), .ZN(
        cell_1000_n41) );
  XOR2_X1 cell_1000_U15 ( .A(cell_1000_g2_0_2_), .B(cell_1000_g2_0_1_), .Z(
        cell_1000_n2) );
  XOR2_X1 cell_1000_U14 ( .A(cell_1000_g5_0_2_), .B(cell_1000_g5_0_1_), .Z(
        cell_1000_n67) );
  XNOR2_X1 cell_1000_U13 ( .A(cell_1000_n1), .B(signal_1257), .ZN(signal_1436)
         );
  XNOR2_X1 cell_1000_U12 ( .A(cell_1000_n109), .B(1'b0), .ZN(cell_1000_n1) );
  XOR2_X1 cell_1000_U11 ( .A(cell_1000_g10_1_2_), .B(cell_1000_g10_1_3_), .Z(
        cell_1000_n109) );
  XNOR2_X1 cell_1000_U10 ( .A(cell_1000_n4), .B(cell_1000_n136), .ZN(
        signal_1472) );
  XNOR2_X1 cell_1000_U9 ( .A(cell_1000_g5_1_2_), .B(cell_1000_g5_1_3_), .ZN(
        cell_1000_n136) );
  XNOR2_X1 cell_1000_U8 ( .A(signal_1245), .B(cell_1000_n7), .ZN(cell_1000_n4)
         );
  XNOR2_X1 cell_1000_U7 ( .A(cell_1000_g2_1_2_), .B(cell_1000_g2_1_3_), .ZN(
        cell_1000_n7) );
  XNOR2_X1 cell_1000_U6 ( .A(cell_1000_n11), .B(cell_1000_n150), .ZN(
        signal_1476) );
  XNOR2_X1 cell_1000_U5 ( .A(cell_1000_g4_1_2_), .B(cell_1000_g4_1_3_), .ZN(
        cell_1000_n150) );
  XNOR2_X1 cell_1000_U4 ( .A(signal_1233), .B(cell_1000_n14), .ZN(
        cell_1000_n11) );
  XNOR2_X1 cell_1000_U3 ( .A(cell_1000_g1_1_2_), .B(cell_1000_g1_1_3_), .ZN(
        cell_1000_n14) );
  XNOR2_X1 cell_1000_U2 ( .A(cell_1000_g4_0_2_), .B(cell_1000_n10), .ZN(
        signal_835) );
  XNOR2_X1 cell_1000_U1 ( .A(cell_1000_g1_0_2_), .B(signal_1143), .ZN(
        cell_1000_n10) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n379), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n377), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n378), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n372), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n368), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n366), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n363), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n360), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n358), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A2(Fresh[3]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313), .A2(Fresh[3]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311), .A2(Fresh[3]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n377), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n373), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A3(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U151 ( .A1(
        Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U138 ( .A1(
        Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n376), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U124 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U118 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U114 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .B(Fresh[2]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A3(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252), .B(Fresh[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U88 ( .B1(
        Ciphertext_s0[48]), .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), 
        .A(Ciphertext_s0[50]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U86 ( .A1(
        Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U84 ( .A1(
        Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U83 ( .A1(Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .A2(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U75 ( .A1(Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n225), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n223), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n221), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U68 ( .A1(
        Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n220), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n219), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n218), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n225), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n217), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U59 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n223), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U55 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A3(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n216), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n224), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n222), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U50 ( .A(Fresh[1]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n215), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n224), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U46 ( .A1(
        Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U42 ( .A1(
        Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n213), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U36 ( .A1(
        Ciphertext_s0[49]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n212), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U28 ( .A1(
        Ciphertext_s0[49]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .A2(Ciphertext_s0[50]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n211), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U17 ( .A1(
        Ciphertext_s0[49]), .A2(Ciphertext_s0[51]), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U13 ( .A(Fresh[0]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U12 ( .A1(Ciphertext_s0[49]), .A2(Ciphertext_s0[48]), .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U11 ( .A(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U10 ( .A(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U7 ( .A(Ciphertext_s0[50]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U6 ( .A(Ciphertext_s0[51]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U1 ( .A(Fresh[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U88 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n68), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n67), .ZN(cell_1000_g0_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U87 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n67) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n68) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53), .ZN(cell_1000_g0_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39), .ZN(cell_1000_g0_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25), .ZN(cell_1000_g0_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U18 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U12 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U7 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U4 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8) );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n83), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n82), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n81), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n80), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n79), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n78), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n77), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n76), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n75), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n74), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n73), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n72), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n71), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n70), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n69), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_0_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[0]), .CK(clk), .Q(cell_1000_GHPC_Gadget_0_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g0_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[1]), .CK(clk), .Q(cell_1000_GHPC_Gadget_0_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g0_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[2]), .CK(clk), .Q(cell_1000_GHPC_Gadget_0_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g0_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[3]), .CK(clk), .Q(cell_1000_GHPC_Gadget_0_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g0_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n379), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n377), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n378), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n372), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n368), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n366), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n363), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n360), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n358), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A2(Fresh[7]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313), .A2(Fresh[7]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311), .A2(Fresh[7]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n377), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n373), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A3(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U151 ( .A1(
        Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U138 ( .A1(
        Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n376), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U124 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U118 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U114 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .B(Fresh[6]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A3(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252), .B(Fresh[5]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U88 ( .B1(
        Ciphertext_s0[52]), .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), 
        .A(Ciphertext_s0[54]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U86 ( .A1(
        Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U84 ( .A1(
        Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U83 ( .A1(Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .A2(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U75 ( .A1(Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n225), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n223), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n221), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U68 ( .A1(
        Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n220), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n219), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n218), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n225), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n217), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U59 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n223), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U55 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A3(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n216), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n224), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n222), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U50 ( .A(Fresh[5]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n215), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n224), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U46 ( .A1(
        Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U42 ( .A1(
        Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n213), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U36 ( .A1(
        Ciphertext_s0[53]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n212), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U28 ( .A1(
        Ciphertext_s0[53]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .A2(Ciphertext_s0[54]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n211), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U17 ( .A1(
        Ciphertext_s0[53]), .A2(Ciphertext_s0[55]), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U13 ( .A(Fresh[4]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U12 ( .A1(Ciphertext_s0[53]), .A2(Ciphertext_s0[52]), .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U11 ( .A(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U10 ( .A(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U7 ( .A(Ciphertext_s0[54]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U6 ( .A(Ciphertext_s0[55]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U1 ( .A(Fresh[7]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n231), .ZN(cell_1000_g1_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n217), .ZN(cell_1000_g1_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n203), .ZN(cell_1000_g1_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189), .ZN(cell_1000_g1_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_1_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[4]), .CK(clk), .Q(cell_1000_GHPC_Gadget_1_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g1_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[5]), .CK(clk), .Q(cell_1000_GHPC_Gadget_1_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g1_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[6]), .CK(clk), .Q(cell_1000_GHPC_Gadget_1_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g1_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[7]), .CK(clk), .Q(cell_1000_GHPC_Gadget_1_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g1_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[59]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[57]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[56]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n379), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n377), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n378), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n372), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n368), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n366), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n363), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n360), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n358), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A2(Fresh[11]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313), .A2(Fresh[11]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311), .A2(Fresh[11]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n377), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n373), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A3(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U151 ( .A1(
        Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U138 ( .A1(
        Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n376), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U124 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U118 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U114 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .B(Fresh[10]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A3(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252), .B(Fresh[9]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U88 ( .B1(
        Ciphertext_s0[56]), .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), 
        .A(Ciphertext_s0[58]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U86 ( .A1(
        Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U84 ( .A1(
        Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U83 ( .A1(Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .A2(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U75 ( .A1(Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n225), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n223), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n221), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U68 ( .A1(
        Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n220), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n219), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n218), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n225), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n217), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U59 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n223), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U55 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A3(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n216), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n224), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n222), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U50 ( .A(Fresh[9]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n215), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n224), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U46 ( .A1(
        Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U42 ( .A1(
        Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n213), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U36 ( .A1(
        Ciphertext_s0[57]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n212), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U28 ( .A1(
        Ciphertext_s0[57]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .A2(Ciphertext_s0[58]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n211), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U17 ( .A1(
        Ciphertext_s0[57]), .A2(Ciphertext_s0[59]), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U13 ( .A(Fresh[8]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U12 ( .A1(Ciphertext_s0[57]), .A2(Ciphertext_s0[56]), .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U11 ( .A(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U10 ( .A(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U7 ( .A(Ciphertext_s0[58]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U6 ( .A(Ciphertext_s0[59]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U1 ( .A(Fresh[11]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n231), .ZN(cell_1000_g2_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n217), .ZN(cell_1000_g2_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n203), .ZN(cell_1000_g2_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189), .ZN(cell_1000_g2_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_2_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[8]), .CK(clk), .Q(cell_1000_GHPC_Gadget_2_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g2_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[9]), .CK(clk), .Q(cell_1000_GHPC_Gadget_2_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g2_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[10]), .CK(clk), .Q(cell_1000_GHPC_Gadget_2_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g2_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[11]), .CK(clk), .Q(cell_1000_GHPC_Gadget_2_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g2_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n379), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n377), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n378), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n372), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n368), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n366), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n363), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n360), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n358), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A2(Fresh[15]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313), .A2(Fresh[15]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311), .A2(Fresh[15]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n377), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n373), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A3(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U151 ( .A1(
        Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U138 ( .A1(
        Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n376), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U124 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U118 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U114 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .B(Fresh[14]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A3(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252), .B(Fresh[13]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U88 ( .B1(
        Ciphertext_s0[24]), .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), 
        .A(Ciphertext_s0[26]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U86 ( .A1(
        Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U84 ( .A1(
        Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U83 ( .A1(Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .A2(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U75 ( .A1(Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n225), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n223), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n221), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U68 ( .A1(
        Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n220), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n219), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n218), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n225), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n217), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U59 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n223), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U55 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A3(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n216), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n224), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n222), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U50 ( .A(Fresh[13]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n215), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n224), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U46 ( .A1(
        Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U42 ( .A1(
        Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n213), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U36 ( .A1(
        Ciphertext_s0[25]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n212), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U28 ( .A1(
        Ciphertext_s0[25]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .A2(Ciphertext_s0[26]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n211), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U17 ( .A1(
        Ciphertext_s0[25]), .A2(Ciphertext_s0[27]), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U13 ( .A(Fresh[12]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U12 ( .A1(Ciphertext_s0[25]), .A2(Ciphertext_s0[24]), .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U11 ( .A(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U10 ( .A(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U7 ( .A(Ciphertext_s0[26]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U6 ( .A(Ciphertext_s0[27]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U1 ( .A(Fresh[15]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n231), .ZN(cell_1000_g3_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n217), .ZN(cell_1000_g3_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n203), .ZN(cell_1000_g3_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189), .ZN(cell_1000_g3_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_3_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[12]), .CK(clk), .Q(cell_1000_GHPC_Gadget_3_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g3_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[13]), .CK(clk), .Q(cell_1000_GHPC_Gadget_3_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g3_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[14]), .CK(clk), .Q(cell_1000_GHPC_Gadget_3_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g3_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[15]), .CK(clk), .Q(cell_1000_GHPC_Gadget_3_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g3_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n379), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n377), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n378), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n372), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n368), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n366), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n363), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n360), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n358), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A2(Fresh[19]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313), .A2(Fresh[19]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311), .A2(Fresh[19]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n377), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n373), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A3(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U151 ( .A1(
        Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U138 ( .A1(
        Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n376), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U124 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U118 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U114 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .B(Fresh[18]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A3(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252), .B(Fresh[17]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U88 ( .B1(
        Ciphertext_s0[28]), .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), 
        .A(Ciphertext_s0[30]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U86 ( .A1(
        Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U84 ( .A1(
        Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U83 ( .A1(Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .A2(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U75 ( .A1(Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n225), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n223), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n221), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U68 ( .A1(
        Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n220), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n219), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n218), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n225), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n217), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U59 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n223), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U55 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A3(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n216), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n224), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n222), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U50 ( .A(Fresh[17]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n215), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n224), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U46 ( .A1(
        Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U42 ( .A1(
        Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n213), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U36 ( .A1(
        Ciphertext_s0[29]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n212), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U28 ( .A1(
        Ciphertext_s0[29]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .A2(Ciphertext_s0[30]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n211), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U17 ( .A1(
        Ciphertext_s0[29]), .A2(Ciphertext_s0[31]), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U13 ( .A(Fresh[16]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U12 ( .A1(Ciphertext_s0[29]), .A2(Ciphertext_s0[28]), .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U11 ( .A(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U10 ( .A(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U7 ( .A(Ciphertext_s0[30]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U6 ( .A(Ciphertext_s0[31]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U1 ( .A(Fresh[19]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n231), .ZN(cell_1000_g4_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n217), .ZN(cell_1000_g4_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n203), .ZN(cell_1000_g4_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189), .ZN(cell_1000_g4_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_4_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[16]), .CK(clk), .Q(cell_1000_GHPC_Gadget_4_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g4_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[17]), .CK(clk), .Q(cell_1000_GHPC_Gadget_4_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g4_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[18]), .CK(clk), .Q(cell_1000_GHPC_Gadget_4_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g4_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[19]), .CK(clk), .Q(cell_1000_GHPC_Gadget_4_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g4_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n379), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n377), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n378), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n372), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n368), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n366), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n363), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n360), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n358), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A2(Fresh[23]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313), .A2(Fresh[23]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311), .A2(Fresh[23]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n377), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n373), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A3(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U151 ( .A1(
        Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U138 ( .A1(
        Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n376), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U124 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U118 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U114 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .B(Fresh[22]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A3(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252), .B(Fresh[21]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U88 ( .B1(
        Ciphertext_s0[16]), .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), 
        .A(Ciphertext_s0[18]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U86 ( .A1(
        Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U84 ( .A1(
        Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U83 ( .A1(Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .A2(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U75 ( .A1(Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n225), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n223), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n221), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U68 ( .A1(
        Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n220), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n219), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n218), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n225), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n217), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U59 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n223), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U55 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A3(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n216), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n224), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n222), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U50 ( .A(Fresh[21]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n215), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n224), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U46 ( .A1(
        Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U42 ( .A1(
        Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n213), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U36 ( .A1(
        Ciphertext_s0[17]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n212), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U28 ( .A1(
        Ciphertext_s0[17]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .A2(Ciphertext_s0[18]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n211), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U17 ( .A1(
        Ciphertext_s0[17]), .A2(Ciphertext_s0[19]), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U13 ( .A(Fresh[20]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U12 ( .A1(Ciphertext_s0[17]), .A2(Ciphertext_s0[16]), .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U11 ( .A(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U10 ( .A(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U7 ( .A(Ciphertext_s0[18]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U6 ( .A(Ciphertext_s0[19]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U1 ( .A(Fresh[23]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n231), .ZN(cell_1000_g5_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n217), .ZN(cell_1000_g5_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n203), .ZN(cell_1000_g5_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189), .ZN(cell_1000_g5_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_5_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[20]), .CK(clk), .Q(cell_1000_GHPC_Gadget_5_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g5_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[21]), .CK(clk), .Q(cell_1000_GHPC_Gadget_5_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g5_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[22]), .CK(clk), .Q(cell_1000_GHPC_Gadget_5_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g5_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[23]), .CK(clk), .Q(cell_1000_GHPC_Gadget_5_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g5_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n379), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n377), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n378), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n372), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n368), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n366), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n363), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n360), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n358), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A2(Fresh[27]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313), .A2(Fresh[27]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311), .A2(Fresh[27]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n377), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n373), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A3(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U151 ( .A1(
        Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U138 ( .A1(
        Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n376), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U124 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U118 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U114 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .B(Fresh[26]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A3(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252), .B(Fresh[25]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U88 ( .B1(
        Ciphertext_s0[36]), .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), 
        .A(Ciphertext_s0[38]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U86 ( .A1(
        Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U84 ( .A1(
        Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U83 ( .A1(Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .A2(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U75 ( .A1(Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n225), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n223), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n221), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U68 ( .A1(
        Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n220), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n219), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n218), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n225), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n217), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U59 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n223), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U55 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A3(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n216), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n224), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n222), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U50 ( .A(Fresh[25]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n215), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n224), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U46 ( .A1(
        Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U42 ( .A1(
        Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n213), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U36 ( .A1(
        Ciphertext_s0[37]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n212), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U28 ( .A1(
        Ciphertext_s0[37]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .A2(Ciphertext_s0[38]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n211), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U17 ( .A1(
        Ciphertext_s0[37]), .A2(Ciphertext_s0[39]), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U13 ( .A(Fresh[24]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U12 ( .A1(Ciphertext_s0[37]), .A2(Ciphertext_s0[36]), .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U11 ( .A(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U10 ( .A(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U7 ( .A(Ciphertext_s0[38]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U6 ( .A(Ciphertext_s0[39]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U1 ( .A(Fresh[27]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n231), .ZN(cell_1000_g6_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n217), .ZN(cell_1000_g6_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n203), .ZN(cell_1000_g6_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189), .ZN(cell_1000_g6_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_6_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[24]), .CK(clk), .Q(cell_1000_GHPC_Gadget_6_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g6_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[25]), .CK(clk), .Q(cell_1000_GHPC_Gadget_6_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g6_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[26]), .CK(clk), .Q(cell_1000_GHPC_Gadget_6_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g6_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[27]), .CK(clk), .Q(cell_1000_GHPC_Gadget_6_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g6_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n379), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n377), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n378), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n372), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n368), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n366), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n363), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n360), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n358), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A2(Fresh[31]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313), .A2(Fresh[31]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311), .A2(Fresh[31]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n377), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n373), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A3(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U151 ( .A1(
        Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U138 ( .A1(
        Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n376), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U124 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U118 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U114 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .B(Fresh[30]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A3(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252), .B(Fresh[29]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U88 ( .B1(
        Ciphertext_s0[40]), .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), 
        .A(Ciphertext_s0[42]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U86 ( .A1(
        Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U84 ( .A1(
        Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U83 ( .A1(Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .A2(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U75 ( .A1(Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n225), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n223), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n221), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U68 ( .A1(
        Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n220), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n219), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n218), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n225), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n217), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U59 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n223), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U55 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A3(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n216), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n224), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n222), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U50 ( .A(Fresh[29]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n215), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n224), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U46 ( .A1(
        Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U42 ( .A1(
        Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n213), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U36 ( .A1(
        Ciphertext_s0[41]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n212), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U28 ( .A1(
        Ciphertext_s0[41]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .A2(Ciphertext_s0[42]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n211), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U17 ( .A1(
        Ciphertext_s0[41]), .A2(Ciphertext_s0[43]), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U13 ( .A(Fresh[28]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U12 ( .A1(Ciphertext_s0[41]), .A2(Ciphertext_s0[40]), .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U11 ( .A(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U10 ( .A(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U7 ( .A(Ciphertext_s0[42]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U6 ( .A(Ciphertext_s0[43]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U1 ( .A(Fresh[31]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n231), .ZN(cell_1000_g7_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n217), .ZN(cell_1000_g7_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n203), .ZN(cell_1000_g7_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189), .ZN(cell_1000_g7_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_7_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[28]), .CK(clk), .Q(cell_1000_GHPC_Gadget_7_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g7_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[29]), .CK(clk), .Q(cell_1000_GHPC_Gadget_7_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g7_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[30]), .CK(clk), .Q(cell_1000_GHPC_Gadget_7_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g7_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[31]), .CK(clk), .Q(cell_1000_GHPC_Gadget_7_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g7_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n379), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n377), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n378), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n372), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n368), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n366), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n363), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n360), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n358), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A2(Fresh[35]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313), .A2(Fresh[35]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311), .A2(Fresh[35]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n377), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n373), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A3(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U151 ( .A1(
        Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U138 ( .A1(
        Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n376), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U124 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U118 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U114 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .B(Fresh[34]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A3(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252), .B(Fresh[33]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U88 ( .B1(
        Ciphertext_s0[20]), .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), 
        .A(Ciphertext_s0[22]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U86 ( .A1(
        Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U84 ( .A1(
        Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U83 ( .A1(Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .A2(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U75 ( .A1(Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n225), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n223), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n221), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U68 ( .A1(
        Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n220), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n219), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n218), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n225), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n217), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U59 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n223), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U55 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A3(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n216), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n224), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n222), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U50 ( .A(Fresh[33]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n215), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n224), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U46 ( .A1(
        Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U42 ( .A1(
        Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n213), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U36 ( .A1(
        Ciphertext_s0[21]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n212), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U28 ( .A1(
        Ciphertext_s0[21]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .A2(Ciphertext_s0[22]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n211), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U17 ( .A1(
        Ciphertext_s0[21]), .A2(Ciphertext_s0[23]), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U13 ( .A(Fresh[32]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U12 ( .A1(Ciphertext_s0[21]), .A2(Ciphertext_s0[20]), .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U11 ( .A(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U10 ( .A(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U7 ( .A(Ciphertext_s0[22]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U6 ( .A(Ciphertext_s0[23]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U1 ( .A(Fresh[35]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n231), .ZN(cell_1000_g8_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n217), .ZN(cell_1000_g8_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n203), .ZN(cell_1000_g8_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189), .ZN(cell_1000_g8_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_8_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[32]), .CK(clk), .Q(cell_1000_GHPC_Gadget_8_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g8_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[33]), .CK(clk), .Q(cell_1000_GHPC_Gadget_8_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g8_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[34]), .CK(clk), .Q(cell_1000_GHPC_Gadget_8_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g8_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[35]), .CK(clk), .Q(cell_1000_GHPC_Gadget_8_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g8_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n379), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n377), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n378), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n372), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n368), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n366), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n363), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n360), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n358), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A2(Fresh[39]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313), .A2(Fresh[39]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311), .A2(Fresh[39]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n377), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n373), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A3(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U151 ( .A1(
        Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U138 ( .A1(
        Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n376), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U124 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U118 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U114 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .B(Fresh[38]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A3(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252), .B(Fresh[37]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U88 ( .B1(
        Ciphertext_s0[32]), .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), 
        .A(Ciphertext_s0[34]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U86 ( .A1(
        Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), 
        .B1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U84 ( .A1(
        Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), 
        .B1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U83 ( .A1(Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .A2(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U75 ( .A1(Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n225), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n223), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n221), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U68 ( .A1(
        Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n220), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n219), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n218), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n225), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n217), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U59 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n223), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U55 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A3(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n216), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n224), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n222), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U50 ( .A(Fresh[37]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n215), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n224), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U46 ( .A1(
        Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U42 ( .A1(
        Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n213), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U36 ( .A1(
        Ciphertext_s0[33]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n212), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U28 ( .A1(
        Ciphertext_s0[33]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .A2(Ciphertext_s0[34]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n211), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U17 ( .A1(
        Ciphertext_s0[33]), .A2(Ciphertext_s0[35]), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U13 ( .A(Fresh[36]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U12 ( .A1(Ciphertext_s0[33]), .A2(Ciphertext_s0[32]), .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275)
         );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U11 ( .A(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U10 ( .A(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U7 ( .A(Ciphertext_s0[34]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U6 ( .A(Ciphertext_s0[35]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U1 ( .A(Fresh[39]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n231), .ZN(cell_1000_g9_1_3_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n217), .ZN(cell_1000_g9_1_2_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n203), .ZN(cell_1000_g9_1_1_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189), .ZN(cell_1000_g9_1_0_)
         );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168) );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[48]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[49]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[50]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[51]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[52]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[53]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[54]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[55]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[56]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[57]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[58]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[59]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[60]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[61]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[62]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_0_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[63]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[32]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[33]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[34]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[35]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[36]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[37]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[38]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[39]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[40]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[41]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[42]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[43]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[44]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[45]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[46]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_1_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[47]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[16]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[17]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[18]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[19]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[20]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[21]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[22]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[23]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[24]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[25]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[26]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[27]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[28]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[29]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[30]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_2_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[31]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_10_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[10]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_11_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[11]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_12_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[12]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_13_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[13]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_14_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[14]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step2_inst_step2_ins_3_15_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_9_inst_Step2_inst_Step2_reg[15]), .QN()
         );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[36]), .CK(clk), .Q(cell_1000_GHPC_Gadget_9_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g9_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[37]), .CK(clk), .Q(cell_1000_GHPC_Gadget_9_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g9_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[38]), .CK(clk), .Q(cell_1000_GHPC_Gadget_9_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g9_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[39]), .CK(clk), .Q(cell_1000_GHPC_Gadget_9_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g9_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[63]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[61]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[60]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n379), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n377), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n378), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n372), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n368), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n366), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n363), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n360), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n358), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A2(Fresh[43]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313), .A2(Fresh[43]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311), .A2(Fresh[43]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n377), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n373), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A3(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U151 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U138 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n376), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U124 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U118 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U114 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .B(Fresh[42]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A3(
        Ciphertext_s0[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252), .B(Fresh[41]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U88 ( .B1(
        Ciphertext_s0[60]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .A(Ciphertext_s0[62]), .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U86 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U84 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U83 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .A2(
        Ciphertext_s0[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U75 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n225), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n223), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n221), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U68 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n220), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n219), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n218), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n225), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n217), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U59 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n223), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U55 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A3(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n216), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n224), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n222), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U50 ( .A(Fresh[41]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n215), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n224), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U46 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U42 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n213), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U36 ( .A1(
        Ciphertext_s0[61]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n212), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U28 ( .A1(
        Ciphertext_s0[61]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .A2(
        Ciphertext_s0[62]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n211), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U17 ( .A1(
        Ciphertext_s0[61]), .A2(Ciphertext_s0[63]), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U13 ( .A(Fresh[40]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U12 ( .A1(
        Ciphertext_s0[61]), .A2(Ciphertext_s0[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U11 ( .A(Ciphertext_s0[61]), .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U10 ( .A(Ciphertext_s0[60]), .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U7 ( .A(Ciphertext_s0[62]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U6 ( .A(Ciphertext_s0[63]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U1 ( .A(Fresh[43]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n231), .ZN(cell_1000_g10_1_3_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n217), .ZN(cell_1000_g10_1_2_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n203), .ZN(cell_1000_g10_1_1_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189), .ZN(cell_1000_g10_1_0_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[40]), .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g10_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[41]), .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g10_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[42]), .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g10_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[43]), .CK(clk), .Q(cell_1000_GHPC_Gadget_10_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g10_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n379), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n377), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n378), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n372), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n368), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n366), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n363), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n360), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n358), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A2(Fresh[47]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313), .A2(Fresh[47]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311), .A2(Fresh[47]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n377), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n373), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A3(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U151 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U138 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n376), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U124 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U118 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U114 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .B(Fresh[46]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A3(
        Ciphertext_s0[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252), .B(Fresh[45]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U88 ( .B1(
        Ciphertext_s0[12]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .A(Ciphertext_s0[14]), .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U86 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U84 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U83 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .A2(
        Ciphertext_s0[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U75 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n225), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n223), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n221), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U68 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n220), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n219), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n218), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n225), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n217), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U59 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n223), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U55 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A3(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n216), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n224), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n222), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U50 ( .A(Fresh[45]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n215), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n224), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U46 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U42 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n213), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U36 ( .A1(
        Ciphertext_s0[13]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n212), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U28 ( .A1(
        Ciphertext_s0[13]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .A2(
        Ciphertext_s0[14]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n211), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U17 ( .A1(
        Ciphertext_s0[13]), .A2(Ciphertext_s0[15]), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U13 ( .A(Fresh[44]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U12 ( .A1(
        Ciphertext_s0[13]), .A2(Ciphertext_s0[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U11 ( .A(Ciphertext_s0[13]), .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U10 ( .A(Ciphertext_s0[12]), .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U7 ( .A(Ciphertext_s0[14]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U6 ( .A(Ciphertext_s0[15]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U1 ( .A(Fresh[47]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n231), .ZN(cell_1000_g11_1_3_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n217), .ZN(cell_1000_g11_1_2_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n203), .ZN(cell_1000_g11_1_1_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189), .ZN(cell_1000_g11_1_0_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173) );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[44]), .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g11_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[45]), .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g11_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[46]), .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g11_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[47]), .CK(clk), .Q(cell_1000_GHPC_Gadget_11_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g11_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n379), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n377), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n378), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n372), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n368), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n366), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n363), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n360), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n358), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A2(Fresh[51]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313), .A2(Fresh[51]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311), .A2(Fresh[51]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n377), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n373), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A3(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U151 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U138 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n376), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U124 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U118 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U114 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .B(Fresh[50]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A3(Ciphertext_s0[0]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252), .B(Fresh[49]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U88 ( .B1(
        Ciphertext_s0[0]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .A(Ciphertext_s0[2]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242)
         );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U86 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U84 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .B1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U83 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .A2(Ciphertext_s0[0]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U75 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n225), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n223), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n221), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U68 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n220), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n219), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n218), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n225), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n217), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U59 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n223), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U55 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A3(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n216), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n224), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n222), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U50 ( .A(Fresh[49]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n215), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n224), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U46 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U42 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n213), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U36 ( .A1(
        Ciphertext_s0[1]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n212), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U28 ( .A1(
        Ciphertext_s0[1]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .A2(Ciphertext_s0[2]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n211), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U17 ( .A1(
        Ciphertext_s0[1]), .A2(Ciphertext_s0[3]), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U13 ( .A(Fresh[48]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U12 ( .A1(
        Ciphertext_s0[1]), .A2(Ciphertext_s0[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U11 ( .A(Ciphertext_s0[1]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U10 ( .A(Ciphertext_s0[0]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U7 ( .A(Ciphertext_s0[2]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U6 ( .A(Ciphertext_s0[3]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U1 ( .A(Fresh[51]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n231), .ZN(cell_1000_g12_1_3_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n217), .ZN(cell_1000_g12_1_2_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n203), .ZN(cell_1000_g12_1_1_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189), .ZN(cell_1000_g12_1_0_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[48]), .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g12_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[49]), .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g12_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[50]), .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g12_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[51]), .CK(clk), .Q(cell_1000_GHPC_Gadget_12_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g12_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n379), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n377), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n378), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n372), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n368), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n366), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n363), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n360), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n358), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A2(Fresh[55]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313), .A2(Fresh[55]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311), .A2(Fresh[55]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n377), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n373), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A3(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U151 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U138 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n376), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U124 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U118 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U114 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .B(Fresh[54]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A3(Ciphertext_s0[4]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252), .B(Fresh[53]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U88 ( .B1(
        Ciphertext_s0[4]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .A(Ciphertext_s0[6]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242)
         );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U86 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U84 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .B1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U83 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .A2(Ciphertext_s0[4]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U75 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n225), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n223), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n221), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U68 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n220), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n219), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n218), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n225), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n217), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U59 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n223), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U55 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A3(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n216), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n224), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n222), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U50 ( .A(Fresh[53]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n215), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n224), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U46 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U42 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n213), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U36 ( .A1(
        Ciphertext_s0[5]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n212), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U28 ( .A1(
        Ciphertext_s0[5]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .A2(Ciphertext_s0[6]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n211), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U17 ( .A1(
        Ciphertext_s0[5]), .A2(Ciphertext_s0[7]), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U13 ( .A(Fresh[52]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U12 ( .A1(
        Ciphertext_s0[5]), .A2(Ciphertext_s0[4]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U11 ( .A(Ciphertext_s0[5]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U10 ( .A(Ciphertext_s0[4]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U7 ( .A(Ciphertext_s0[6]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U6 ( .A(Ciphertext_s0[7]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U1 ( .A(Fresh[55]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n231), .ZN(cell_1000_g13_1_3_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n217), .ZN(cell_1000_g13_1_2_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n203), .ZN(cell_1000_g13_1_1_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189), .ZN(cell_1000_g13_1_0_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173) );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[52]), .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g13_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[53]), .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g13_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[54]), .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g13_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[55]), .CK(clk), .Q(cell_1000_GHPC_Gadget_13_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g13_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n379), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n377), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n378), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n372), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n368), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n366), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n363), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n360), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n358), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A2(Fresh[59]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313), .A2(Fresh[59]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311), .A2(Fresh[59]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n377), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n373), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A3(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U151 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U138 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n376), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U124 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U118 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U114 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .B(Fresh[58]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A3(
        Ciphertext_s0[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252), .B(Fresh[57]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U88 ( .B1(
        Ciphertext_s0[44]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .A(Ciphertext_s0[46]), .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U86 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U84 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U83 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .A2(
        Ciphertext_s0[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U75 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n225), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n223), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n221), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U68 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n220), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n219), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n218), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n225), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n217), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U59 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n223), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U55 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A3(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n216), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n224), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n222), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U50 ( .A(Fresh[57]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n215), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n224), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U46 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U42 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n213), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U36 ( .A1(
        Ciphertext_s0[45]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n212), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U28 ( .A1(
        Ciphertext_s0[45]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .A2(
        Ciphertext_s0[46]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n211), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U17 ( .A1(
        Ciphertext_s0[45]), .A2(Ciphertext_s0[47]), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U13 ( .A(Fresh[56]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U12 ( .A1(
        Ciphertext_s0[45]), .A2(Ciphertext_s0[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U11 ( .A(Ciphertext_s0[45]), .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U10 ( .A(Ciphertext_s0[44]), .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U7 ( .A(Ciphertext_s0[46]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U6 ( .A(Ciphertext_s0[47]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U1 ( .A(Fresh[59]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n231), .ZN(cell_1000_g14_1_3_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n217), .ZN(cell_1000_g14_1_2_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n203), .ZN(cell_1000_g14_1_1_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189), .ZN(cell_1000_g14_1_0_) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[56]), .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g14_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[57]), .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g14_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[58]), .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g14_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[59]), .CK(clk), .Q(cell_1000_GHPC_Gadget_14_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g14_0_3_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U226 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n379), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n378), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n176) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U225 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n377), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n379) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U224 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n378), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n375), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[8]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U223 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n373), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n375) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U222 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n372), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n378) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U221 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n368), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[7]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U220 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n366), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n365), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n368) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U219 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n365) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U218 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n363), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n367), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[6]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U217 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n367) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U216 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n360), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n363) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U215 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n358), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[5]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U214 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n358) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U213 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U212 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U211 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U210 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[3]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U209 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U208 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U207 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A2(Fresh[63]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U206 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U205 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U204 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[1]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U203 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n376), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U202 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U201 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U200 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[13]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U199 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U198 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U197 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[12]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U195 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[11]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U192 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U190 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[9]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U188 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U187 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U184 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313), .A2(Fresh[63]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U183 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n370) );
  OAI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311), .A2(Fresh[63]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n371) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U181 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U180 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[24]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n377), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U178 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n377) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U177 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[23]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U176 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n373), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U175 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n373) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U174 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n366), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[22]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n366) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U172 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U171 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n360), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U170 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n360) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U169 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U168 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[20]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U166 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U164 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[19]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U163 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U162 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350) );
  NOR3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U161 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A3(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U160 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U159 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[18]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U158 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U157 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U156 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[17]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U155 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U154 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U153 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U152 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U151 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U150 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[16]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U149 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[30]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[29]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U141 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U138 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[28]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U136 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n376), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n376) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U134 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U132 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[27]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U130 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U129 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U128 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U126 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U125 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U124 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[25]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U122 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U121 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U119 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U118 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U117 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[15]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U116 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U114 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U113 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U112 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .B(Fresh[62]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U109 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[40]) );
  OAI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U107 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U106 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[39]) );
  OAI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U104 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n372), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n369) );
  NOR3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U103 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A3(Ciphertext_s0[8]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n372) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U102 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U101 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252), .B(Fresh[61]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U100 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[38]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U97 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U96 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n361) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U94 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n362) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U93 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[36]) );
  OAI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U92 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[35]) );
  OAI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U89 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U88 ( .B1(
        Ciphertext_s0[8]), .B2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .A(Ciphertext_s0[10]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242)
         );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[34]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U86 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B1(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[33]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U84 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .B1(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U83 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[32]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U81 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U80 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .A2(Ciphertext_s0[8]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U79 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[46]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U78 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U77 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[45]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U75 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[44]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U73 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n225), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n224), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U71 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n223), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U70 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n221), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[43]) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U68 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n220), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n221) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n219), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n218), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U64 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n222), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n225), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n219) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U62 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n225) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U61 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n217), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[41]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U59 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n217) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U57 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U56 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n223), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U55 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238) );
  NAND3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A3(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U53 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n216), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n220), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U52 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n224), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n220) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U51 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n222), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U50 ( .A(Fresh[61]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n215), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n223) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U49 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n224), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n218), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n215) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U48 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n218) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U47 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U46 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n224) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U45 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n216) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U44 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U43 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U42 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n15), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n180) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U40 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n213), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n213) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U38 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U36 ( .A1(
        Ciphertext_s0[9]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U35 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n14), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n212), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n212) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U32 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U31 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n374) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U30 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U28 ( .A1(
        Ciphertext_s0[9]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U27 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .A2(
        Ciphertext_s0[10]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n13), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n211), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n13) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U24 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n211) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U23 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n364) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U21 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n12), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n178) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n210), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n12) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n210) );
  NAND3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U17 ( .A1(
        Ciphertext_s0[9]), .A2(Ciphertext_s0[11]), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n359) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U14 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U13 ( .A(Fresh[60]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n214) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U12 ( .A1(
        Ciphertext_s0[9]), .A2(Ciphertext_s0[8]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U11 ( .A(Ciphertext_s0[9]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U10 ( .A(Ciphertext_s0[8]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U9 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U8 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U7 ( .A(Ciphertext_s0[10]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U6 ( .A(Ciphertext_s0[11]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n223), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n222) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U4 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U1 ( .A(Fresh[63]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n14), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n15), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n13), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n12), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n180), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n179), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n178), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n177), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n176), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[15]), .QN() );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U86 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n232), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n231), .ZN(cell_1000_g15_1[3]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U85 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n230), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n229), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n231) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U84 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n228), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n227), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U83 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n226), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n225), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U82 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[1]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n225) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U81 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[0]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[3]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n226) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U80 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n224), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n223), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n228) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U79 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[12]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n223) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U78 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[10]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[11]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n224) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U77 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n222), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n221), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n230) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U76 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[14]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n221) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U75 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[9]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[8]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n222) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U74 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n220), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n219), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n232) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U73 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[6]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n219) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U72 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[4]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[5]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n220) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U71 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n218), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n217), .ZN(cell_1000_g15_1[2]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U70 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n216), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n215), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n217) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U69 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n214), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n213), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n215) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U68 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n212), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n211), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n213) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U67 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[17]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n211) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U66 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[16]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[19]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n212) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U65 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n210), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n209), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n214) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U64 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[28]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n209) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U63 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[26]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[27]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n210) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U62 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n208), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n207), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n216) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U61 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[30]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n207) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U60 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[25]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[24]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n208) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U59 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n206), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n205), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n218) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[22]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n205) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U57 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[20]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[21]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n206) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U56 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n204), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n203), .ZN(cell_1000_g15_1[1]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U55 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n202), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n201), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n203) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U54 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n201) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U52 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[33]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U51 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[32]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[35]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U50 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U49 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[44]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U48 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[42]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[43]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U47 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n202) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U46 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[46]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U45 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[41]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[40]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U44 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n204) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U43 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[38]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U42 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[36]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[37]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U41 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189), .ZN(cell_1000_g15_1[0]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U40 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U39 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U38 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U37 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[49]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U36 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[48]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[51]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U34 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[60]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U33 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[58]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[59]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U32 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U31 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[62]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U30 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[57]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[56]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U29 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U28 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[54]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U27 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[52]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[53]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U14 ( .A(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U9 ( .A(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171) );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[48]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[49]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[49]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[50]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[51]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[51]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[52]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[53]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[53]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[54]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[55]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[55]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[56]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[57]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[57]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[58]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[59]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[59]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[60]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[61]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[61]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[62]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[63]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_0_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[63]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[32]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[33]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[33]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[34]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[35]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[35]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[36]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[37]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[37]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[38]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[39]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[39]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[40]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[41]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[41]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[42]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[43]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[43]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[44]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[45]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[45]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[46]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[47]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_1_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[47]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[16]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[17]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[17]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[18]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[19]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[19]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[20]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[21]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[21]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[22]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[23]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[23]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[24]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[25]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[25]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[26]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[27]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[27]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[28]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[29]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[29]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[30]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[31]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_2_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[31]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_0_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n84), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_0_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_0_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_0_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[0]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_1_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n85), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_1_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_1_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_1_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[1]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_2_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n86), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_2_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_2_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_2_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[2]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_3_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n87), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_3_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_3_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_3_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[3]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_4_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n88), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_4_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_4_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_4_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[4]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_5_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n89), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[5]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_5_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_5_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_5_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[5]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_6_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n90), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_6_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_6_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_6_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[6]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_7_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n91), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[7]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_7_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_7_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_7_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[7]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_8_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n92), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_8_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_8_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_8_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[8]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_9_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n93), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[9]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_9_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_9_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_9_value), .CK(
        clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[9]), .QN()
         );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_10_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n94), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_10_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_10_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_10_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[10]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_11_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n95), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[11]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_11_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_11_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_11_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[11]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_12_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n96), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_12_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_12_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_12_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[12]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_13_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n97), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[13]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_13_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_13_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_13_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[13]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_14_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n98), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_14_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_14_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_14_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[14]), 
        .QN() );
  AND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_15_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_N122), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[15]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_15_value) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_15_output_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step2_inst_step2_ins_3_15_value), 
        .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_Step2_inst_Step2_reg[15]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins1_0_s_current_state_reg ( 
        .D(Fresh[60]), .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_out0_mid[0]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g15_0[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins1_1_s_current_state_reg ( 
        .D(Fresh[61]), .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_out0_mid[1]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g15_0[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins1_2_s_current_state_reg ( 
        .D(Fresh[62]), .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_out0_mid[2]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g15_0[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins1_3_s_current_state_reg ( 
        .D(Fresh[63]), .CK(clk), .Q(cell_1000_GHPC_Gadget_15_inst_out0_mid[3]), 
        .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g15_0[3]), .QN() );
  DFF_X1 cell_65_s_reg_0_s_current_state_reg ( .D(signal_840), .CK(signal_1676), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 cell_65_s_reg_1_s_current_state_reg ( .D(signal_1611), .CK(
        signal_1676), .Q(Ciphertext_s1[63]), .QN() );
  DFF_X1 cell_67_s_reg_0_s_current_state_reg ( .D(signal_841), .CK(signal_1676), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 cell_67_s_reg_1_s_current_state_reg ( .D(signal_1609), .CK(
        signal_1676), .Q(Ciphertext_s1[62]), .QN() );
  DFF_X1 cell_69_s_reg_0_s_current_state_reg ( .D(signal_842), .CK(signal_1676), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 cell_69_s_reg_1_s_current_state_reg ( .D(signal_1607), .CK(
        signal_1676), .Q(Ciphertext_s1[61]), .QN() );
  DFF_X1 cell_71_s_reg_0_s_current_state_reg ( .D(signal_843), .CK(signal_1676), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 cell_71_s_reg_1_s_current_state_reg ( .D(signal_1605), .CK(
        signal_1676), .Q(Ciphertext_s1[60]), .QN() );
  DFF_X1 cell_73_s_reg_0_s_current_state_reg ( .D(signal_844), .CK(signal_1676), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 cell_73_s_reg_1_s_current_state_reg ( .D(signal_1603), .CK(
        signal_1676), .Q(Ciphertext_s1[59]), .QN() );
  DFF_X1 cell_75_s_reg_0_s_current_state_reg ( .D(signal_845), .CK(signal_1676), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 cell_75_s_reg_1_s_current_state_reg ( .D(signal_1601), .CK(
        signal_1676), .Q(Ciphertext_s1[58]), .QN() );
  DFF_X1 cell_77_s_reg_0_s_current_state_reg ( .D(signal_846), .CK(signal_1676), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 cell_77_s_reg_1_s_current_state_reg ( .D(signal_1599), .CK(
        signal_1676), .Q(Ciphertext_s1[57]), .QN() );
  DFF_X1 cell_79_s_reg_0_s_current_state_reg ( .D(signal_847), .CK(signal_1676), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 cell_79_s_reg_1_s_current_state_reg ( .D(signal_1597), .CK(
        signal_1676), .Q(Ciphertext_s1[56]), .QN() );
  DFF_X1 cell_81_s_reg_0_s_current_state_reg ( .D(signal_848), .CK(signal_1676), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 cell_81_s_reg_1_s_current_state_reg ( .D(signal_1595), .CK(
        signal_1676), .Q(Ciphertext_s1[55]), .QN() );
  DFF_X1 cell_83_s_reg_0_s_current_state_reg ( .D(signal_849), .CK(signal_1676), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 cell_83_s_reg_1_s_current_state_reg ( .D(signal_1593), .CK(
        signal_1676), .Q(Ciphertext_s1[54]), .QN() );
  DFF_X1 cell_85_s_reg_0_s_current_state_reg ( .D(signal_850), .CK(signal_1676), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 cell_85_s_reg_1_s_current_state_reg ( .D(signal_1591), .CK(
        signal_1676), .Q(Ciphertext_s1[53]), .QN() );
  DFF_X1 cell_87_s_reg_0_s_current_state_reg ( .D(signal_851), .CK(signal_1676), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 cell_87_s_reg_1_s_current_state_reg ( .D(signal_1589), .CK(
        signal_1676), .Q(Ciphertext_s1[52]), .QN() );
  DFF_X1 cell_89_s_reg_0_s_current_state_reg ( .D(signal_852), .CK(signal_1676), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 cell_89_s_reg_1_s_current_state_reg ( .D(signal_1587), .CK(
        signal_1676), .Q(Ciphertext_s1[51]), .QN() );
  DFF_X1 cell_91_s_reg_0_s_current_state_reg ( .D(signal_853), .CK(signal_1676), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 cell_91_s_reg_1_s_current_state_reg ( .D(signal_1585), .CK(
        signal_1676), .Q(Ciphertext_s1[50]), .QN() );
  DFF_X1 cell_93_s_reg_0_s_current_state_reg ( .D(signal_854), .CK(signal_1676), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 cell_93_s_reg_1_s_current_state_reg ( .D(signal_1583), .CK(
        signal_1676), .Q(Ciphertext_s1[49]), .QN() );
  DFF_X1 cell_95_s_reg_0_s_current_state_reg ( .D(signal_855), .CK(signal_1676), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 cell_95_s_reg_1_s_current_state_reg ( .D(signal_1581), .CK(
        signal_1676), .Q(Ciphertext_s1[48]), .QN() );
  DFF_X1 cell_97_s_reg_0_s_current_state_reg ( .D(signal_856), .CK(signal_1676), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 cell_97_s_reg_1_s_current_state_reg ( .D(signal_1579), .CK(
        signal_1676), .Q(Ciphertext_s1[47]), .QN() );
  DFF_X1 cell_99_s_reg_0_s_current_state_reg ( .D(signal_857), .CK(signal_1676), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 cell_99_s_reg_1_s_current_state_reg ( .D(signal_1577), .CK(
        signal_1676), .Q(Ciphertext_s1[46]), .QN() );
  DFF_X1 cell_101_s_reg_0_s_current_state_reg ( .D(signal_858), .CK(
        signal_1676), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 cell_101_s_reg_1_s_current_state_reg ( .D(signal_1575), .CK(
        signal_1676), .Q(Ciphertext_s1[45]), .QN() );
  DFF_X1 cell_103_s_reg_0_s_current_state_reg ( .D(signal_859), .CK(
        signal_1676), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 cell_103_s_reg_1_s_current_state_reg ( .D(signal_1573), .CK(
        signal_1676), .Q(Ciphertext_s1[44]), .QN() );
  DFF_X1 cell_105_s_reg_0_s_current_state_reg ( .D(signal_860), .CK(
        signal_1676), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 cell_105_s_reg_1_s_current_state_reg ( .D(signal_1571), .CK(
        signal_1676), .Q(Ciphertext_s1[43]), .QN() );
  DFF_X1 cell_107_s_reg_0_s_current_state_reg ( .D(signal_861), .CK(
        signal_1676), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 cell_107_s_reg_1_s_current_state_reg ( .D(signal_1569), .CK(
        signal_1676), .Q(Ciphertext_s1[42]), .QN() );
  DFF_X1 cell_109_s_reg_0_s_current_state_reg ( .D(signal_862), .CK(
        signal_1676), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 cell_109_s_reg_1_s_current_state_reg ( .D(signal_1567), .CK(
        signal_1676), .Q(Ciphertext_s1[41]), .QN() );
  DFF_X1 cell_111_s_reg_0_s_current_state_reg ( .D(signal_863), .CK(
        signal_1676), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 cell_111_s_reg_1_s_current_state_reg ( .D(signal_1565), .CK(
        signal_1676), .Q(Ciphertext_s1[40]), .QN() );
  DFF_X1 cell_113_s_reg_0_s_current_state_reg ( .D(signal_864), .CK(
        signal_1676), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 cell_113_s_reg_1_s_current_state_reg ( .D(signal_1563), .CK(
        signal_1676), .Q(Ciphertext_s1[39]), .QN() );
  DFF_X1 cell_115_s_reg_0_s_current_state_reg ( .D(signal_865), .CK(
        signal_1676), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 cell_115_s_reg_1_s_current_state_reg ( .D(signal_1561), .CK(
        signal_1676), .Q(Ciphertext_s1[38]), .QN() );
  DFF_X1 cell_117_s_reg_0_s_current_state_reg ( .D(signal_866), .CK(
        signal_1676), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 cell_117_s_reg_1_s_current_state_reg ( .D(signal_1559), .CK(
        signal_1676), .Q(Ciphertext_s1[37]), .QN() );
  DFF_X1 cell_119_s_reg_0_s_current_state_reg ( .D(signal_867), .CK(
        signal_1676), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 cell_119_s_reg_1_s_current_state_reg ( .D(signal_1557), .CK(
        signal_1676), .Q(Ciphertext_s1[36]), .QN() );
  DFF_X1 cell_121_s_reg_0_s_current_state_reg ( .D(signal_868), .CK(
        signal_1676), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 cell_121_s_reg_1_s_current_state_reg ( .D(signal_1555), .CK(
        signal_1676), .Q(Ciphertext_s1[35]), .QN() );
  DFF_X1 cell_123_s_reg_0_s_current_state_reg ( .D(signal_869), .CK(
        signal_1676), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 cell_123_s_reg_1_s_current_state_reg ( .D(signal_1553), .CK(
        signal_1676), .Q(Ciphertext_s1[34]), .QN() );
  DFF_X1 cell_125_s_reg_0_s_current_state_reg ( .D(signal_870), .CK(
        signal_1676), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 cell_125_s_reg_1_s_current_state_reg ( .D(signal_1551), .CK(
        signal_1676), .Q(Ciphertext_s1[33]), .QN() );
  DFF_X1 cell_127_s_reg_0_s_current_state_reg ( .D(signal_871), .CK(
        signal_1676), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 cell_127_s_reg_1_s_current_state_reg ( .D(signal_1549), .CK(
        signal_1676), .Q(Ciphertext_s1[32]), .QN() );
  DFF_X1 cell_129_s_reg_0_s_current_state_reg ( .D(signal_872), .CK(
        signal_1676), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 cell_129_s_reg_1_s_current_state_reg ( .D(signal_1547), .CK(
        signal_1676), .Q(Ciphertext_s1[31]), .QN() );
  DFF_X1 cell_131_s_reg_0_s_current_state_reg ( .D(signal_873), .CK(
        signal_1676), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 cell_131_s_reg_1_s_current_state_reg ( .D(signal_1545), .CK(
        signal_1676), .Q(Ciphertext_s1[30]), .QN() );
  DFF_X1 cell_133_s_reg_0_s_current_state_reg ( .D(signal_874), .CK(
        signal_1676), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 cell_133_s_reg_1_s_current_state_reg ( .D(signal_1543), .CK(
        signal_1676), .Q(Ciphertext_s1[29]), .QN() );
  DFF_X1 cell_135_s_reg_0_s_current_state_reg ( .D(signal_875), .CK(
        signal_1676), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 cell_135_s_reg_1_s_current_state_reg ( .D(signal_1541), .CK(
        signal_1676), .Q(Ciphertext_s1[28]), .QN() );
  DFF_X1 cell_137_s_reg_0_s_current_state_reg ( .D(signal_876), .CK(
        signal_1676), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 cell_137_s_reg_1_s_current_state_reg ( .D(signal_1539), .CK(
        signal_1676), .Q(Ciphertext_s1[27]), .QN() );
  DFF_X1 cell_139_s_reg_0_s_current_state_reg ( .D(signal_877), .CK(
        signal_1676), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 cell_139_s_reg_1_s_current_state_reg ( .D(signal_1537), .CK(
        signal_1676), .Q(Ciphertext_s1[26]), .QN() );
  DFF_X1 cell_141_s_reg_0_s_current_state_reg ( .D(signal_878), .CK(
        signal_1676), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 cell_141_s_reg_1_s_current_state_reg ( .D(signal_1535), .CK(
        signal_1676), .Q(Ciphertext_s1[25]), .QN() );
  DFF_X1 cell_143_s_reg_0_s_current_state_reg ( .D(signal_879), .CK(
        signal_1676), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 cell_143_s_reg_1_s_current_state_reg ( .D(signal_1533), .CK(
        signal_1676), .Q(Ciphertext_s1[24]), .QN() );
  DFF_X1 cell_145_s_reg_0_s_current_state_reg ( .D(signal_880), .CK(
        signal_1676), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 cell_145_s_reg_1_s_current_state_reg ( .D(signal_1531), .CK(
        signal_1676), .Q(Ciphertext_s1[23]), .QN() );
  DFF_X1 cell_147_s_reg_0_s_current_state_reg ( .D(signal_881), .CK(
        signal_1676), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 cell_147_s_reg_1_s_current_state_reg ( .D(signal_1529), .CK(
        signal_1676), .Q(Ciphertext_s1[22]), .QN() );
  DFF_X1 cell_149_s_reg_0_s_current_state_reg ( .D(signal_882), .CK(
        signal_1676), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 cell_149_s_reg_1_s_current_state_reg ( .D(signal_1527), .CK(
        signal_1676), .Q(Ciphertext_s1[21]), .QN() );
  DFF_X1 cell_151_s_reg_0_s_current_state_reg ( .D(signal_883), .CK(
        signal_1676), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 cell_151_s_reg_1_s_current_state_reg ( .D(signal_1525), .CK(
        signal_1676), .Q(Ciphertext_s1[20]), .QN() );
  DFF_X1 cell_153_s_reg_0_s_current_state_reg ( .D(signal_884), .CK(
        signal_1676), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 cell_153_s_reg_1_s_current_state_reg ( .D(signal_1523), .CK(
        signal_1676), .Q(Ciphertext_s1[19]), .QN() );
  DFF_X1 cell_155_s_reg_0_s_current_state_reg ( .D(signal_885), .CK(
        signal_1676), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 cell_155_s_reg_1_s_current_state_reg ( .D(signal_1521), .CK(
        signal_1676), .Q(Ciphertext_s1[18]), .QN() );
  DFF_X1 cell_157_s_reg_0_s_current_state_reg ( .D(signal_886), .CK(
        signal_1676), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 cell_157_s_reg_1_s_current_state_reg ( .D(signal_1519), .CK(
        signal_1676), .Q(Ciphertext_s1[17]), .QN() );
  DFF_X1 cell_159_s_reg_0_s_current_state_reg ( .D(signal_887), .CK(
        signal_1676), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 cell_159_s_reg_1_s_current_state_reg ( .D(signal_1517), .CK(
        signal_1676), .Q(Ciphertext_s1[16]), .QN() );
  DFF_X1 cell_161_s_reg_0_s_current_state_reg ( .D(signal_888), .CK(
        signal_1676), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 cell_161_s_reg_1_s_current_state_reg ( .D(signal_1515), .CK(
        signal_1676), .Q(Ciphertext_s1[15]), .QN() );
  DFF_X1 cell_163_s_reg_0_s_current_state_reg ( .D(signal_889), .CK(
        signal_1676), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 cell_163_s_reg_1_s_current_state_reg ( .D(signal_1513), .CK(
        signal_1676), .Q(Ciphertext_s1[14]), .QN() );
  DFF_X1 cell_165_s_reg_0_s_current_state_reg ( .D(signal_890), .CK(
        signal_1676), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 cell_165_s_reg_1_s_current_state_reg ( .D(signal_1511), .CK(
        signal_1676), .Q(Ciphertext_s1[13]), .QN() );
  DFF_X1 cell_167_s_reg_0_s_current_state_reg ( .D(signal_891), .CK(
        signal_1676), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 cell_167_s_reg_1_s_current_state_reg ( .D(signal_1509), .CK(
        signal_1676), .Q(Ciphertext_s1[12]), .QN() );
  DFF_X1 cell_169_s_reg_0_s_current_state_reg ( .D(signal_892), .CK(
        signal_1676), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 cell_169_s_reg_1_s_current_state_reg ( .D(signal_1507), .CK(
        signal_1676), .Q(Ciphertext_s1[11]), .QN() );
  DFF_X1 cell_171_s_reg_0_s_current_state_reg ( .D(signal_893), .CK(
        signal_1676), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 cell_171_s_reg_1_s_current_state_reg ( .D(signal_1505), .CK(
        signal_1676), .Q(Ciphertext_s1[10]), .QN() );
  DFF_X1 cell_173_s_reg_0_s_current_state_reg ( .D(signal_894), .CK(
        signal_1676), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 cell_173_s_reg_1_s_current_state_reg ( .D(signal_1503), .CK(
        signal_1676), .Q(Ciphertext_s1[9]), .QN() );
  DFF_X1 cell_175_s_reg_0_s_current_state_reg ( .D(signal_895), .CK(
        signal_1676), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 cell_175_s_reg_1_s_current_state_reg ( .D(signal_1501), .CK(
        signal_1676), .Q(Ciphertext_s1[8]), .QN() );
  DFF_X1 cell_177_s_reg_0_s_current_state_reg ( .D(signal_896), .CK(
        signal_1676), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 cell_177_s_reg_1_s_current_state_reg ( .D(signal_1499), .CK(
        signal_1676), .Q(Ciphertext_s1[7]), .QN() );
  DFF_X1 cell_179_s_reg_0_s_current_state_reg ( .D(signal_897), .CK(
        signal_1676), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 cell_179_s_reg_1_s_current_state_reg ( .D(signal_1497), .CK(
        signal_1676), .Q(Ciphertext_s1[6]), .QN() );
  DFF_X1 cell_181_s_reg_0_s_current_state_reg ( .D(signal_898), .CK(
        signal_1676), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 cell_181_s_reg_1_s_current_state_reg ( .D(signal_1495), .CK(
        signal_1676), .Q(Ciphertext_s1[5]), .QN() );
  DFF_X1 cell_183_s_reg_0_s_current_state_reg ( .D(signal_899), .CK(
        signal_1676), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 cell_183_s_reg_1_s_current_state_reg ( .D(signal_1493), .CK(
        signal_1676), .Q(Ciphertext_s1[4]), .QN() );
  DFF_X1 cell_185_s_reg_0_s_current_state_reg ( .D(signal_900), .CK(
        signal_1676), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 cell_185_s_reg_1_s_current_state_reg ( .D(signal_1491), .CK(
        signal_1676), .Q(Ciphertext_s1[3]), .QN() );
  DFF_X1 cell_187_s_reg_0_s_current_state_reg ( .D(signal_901), .CK(
        signal_1676), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 cell_187_s_reg_1_s_current_state_reg ( .D(signal_1489), .CK(
        signal_1676), .Q(Ciphertext_s1[2]), .QN() );
  DFF_X1 cell_189_s_reg_0_s_current_state_reg ( .D(signal_902), .CK(
        signal_1676), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 cell_189_s_reg_1_s_current_state_reg ( .D(signal_1487), .CK(
        signal_1676), .Q(Ciphertext_s1[1]), .QN() );
  DFF_X1 cell_191_s_reg_0_s_current_state_reg ( .D(signal_903), .CK(
        signal_1676), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 cell_191_s_reg_1_s_current_state_reg ( .D(signal_1485), .CK(
        signal_1676), .Q(Ciphertext_s1[0]), .QN() );
  DFF_X1 cell_834_s_reg_0_s_current_state_reg ( .D(signal_1036), .CK(
        signal_1676), .Q(signal_1132), .QN() );
  DFF_X1 cell_834_s_reg_1_s_current_state_reg ( .D(signal_1355), .CK(
        signal_1676), .Q(signal_1257), .QN() );
  DFF_X1 cell_836_s_reg_0_s_current_state_reg ( .D(signal_1037), .CK(
        signal_1676), .Q(signal_1133), .QN() );
  DFF_X1 cell_836_s_reg_1_s_current_state_reg ( .D(signal_1352), .CK(
        signal_1676), .Q(signal_1254), .QN() );
  DFF_X1 cell_838_s_reg_0_s_current_state_reg ( .D(signal_1038), .CK(
        signal_1676), .Q(signal_1134), .QN() );
  DFF_X1 cell_838_s_reg_1_s_current_state_reg ( .D(signal_1349), .CK(
        signal_1676), .Q(signal_1251), .QN() );
  DFF_X1 cell_840_s_reg_0_s_current_state_reg ( .D(signal_1039), .CK(
        signal_1676), .Q(signal_1135), .QN() );
  DFF_X1 cell_840_s_reg_1_s_current_state_reg ( .D(signal_1346), .CK(
        signal_1676), .Q(signal_1248), .QN() );
  DFF_X1 cell_842_s_reg_0_s_current_state_reg ( .D(signal_1040), .CK(
        signal_1676), .Q(signal_1136), .QN() );
  DFF_X1 cell_842_s_reg_1_s_current_state_reg ( .D(signal_1343), .CK(
        signal_1676), .Q(signal_1245), .QN() );
  DFF_X1 cell_844_s_reg_0_s_current_state_reg ( .D(signal_1041), .CK(
        signal_1676), .Q(signal_1137), .QN() );
  DFF_X1 cell_844_s_reg_1_s_current_state_reg ( .D(signal_1340), .CK(
        signal_1676), .Q(signal_1242), .QN() );
  DFF_X1 cell_846_s_reg_0_s_current_state_reg ( .D(signal_1042), .CK(
        signal_1676), .Q(signal_1138), .QN() );
  DFF_X1 cell_846_s_reg_1_s_current_state_reg ( .D(signal_1337), .CK(
        signal_1676), .Q(signal_1239), .QN() );
  DFF_X1 cell_848_s_reg_0_s_current_state_reg ( .D(signal_1043), .CK(
        signal_1676), .Q(signal_1139), .QN() );
  DFF_X1 cell_848_s_reg_1_s_current_state_reg ( .D(signal_1334), .CK(
        signal_1676), .Q(signal_1236), .QN() );
  DFF_X1 cell_850_s_reg_0_s_current_state_reg ( .D(signal_1044), .CK(
        signal_1676), .Q(signal_1140), .QN() );
  DFF_X1 cell_850_s_reg_1_s_current_state_reg ( .D(signal_1331), .CK(
        signal_1676), .Q(signal_1233), .QN() );
  DFF_X1 cell_852_s_reg_0_s_current_state_reg ( .D(signal_1045), .CK(
        signal_1676), .Q(signal_1141), .QN() );
  DFF_X1 cell_852_s_reg_1_s_current_state_reg ( .D(signal_1328), .CK(
        signal_1676), .Q(signal_1230), .QN() );
  DFF_X1 cell_854_s_reg_0_s_current_state_reg ( .D(signal_1046), .CK(
        signal_1676), .Q(signal_1142), .QN() );
  DFF_X1 cell_854_s_reg_1_s_current_state_reg ( .D(signal_1325), .CK(
        signal_1676), .Q(signal_1227), .QN() );
  DFF_X1 cell_856_s_reg_0_s_current_state_reg ( .D(signal_1047), .CK(
        signal_1676), .Q(signal_1143), .QN() );
  DFF_X1 cell_856_s_reg_1_s_current_state_reg ( .D(signal_1322), .CK(
        signal_1676), .Q(signal_1224), .QN() );
  DFF_X1 cell_858_s_reg_0_s_current_state_reg ( .D(signal_1048), .CK(
        signal_1676), .Q(signal_1144), .QN() );
  DFF_X1 cell_858_s_reg_1_s_current_state_reg ( .D(signal_1319), .CK(
        signal_1676), .Q(signal_1221), .QN() );
  DFF_X1 cell_860_s_reg_0_s_current_state_reg ( .D(signal_1049), .CK(
        signal_1676), .Q(signal_1145), .QN() );
  DFF_X1 cell_860_s_reg_1_s_current_state_reg ( .D(signal_1316), .CK(
        signal_1676), .Q(signal_1218), .QN() );
  DFF_X1 cell_862_s_reg_0_s_current_state_reg ( .D(signal_1050), .CK(
        signal_1676), .Q(signal_1146), .QN() );
  DFF_X1 cell_862_s_reg_1_s_current_state_reg ( .D(signal_1313), .CK(
        signal_1676), .Q(signal_1215), .QN() );
  DFF_X1 cell_864_s_reg_0_s_current_state_reg ( .D(signal_1051), .CK(
        signal_1676), .Q(signal_1147), .QN() );
  DFF_X1 cell_864_s_reg_1_s_current_state_reg ( .D(signal_1310), .CK(
        signal_1676), .Q(signal_1212), .QN() );
  DFF_X1 cell_866_s_reg_0_s_current_state_reg ( .D(signal_1052), .CK(
        signal_1676), .Q(signal_1148), .QN() );
  DFF_X1 cell_866_s_reg_1_s_current_state_reg ( .D(signal_1307), .CK(
        signal_1676), .Q(signal_1209), .QN() );
  DFF_X1 cell_868_s_reg_0_s_current_state_reg ( .D(signal_1053), .CK(
        signal_1676), .Q(signal_1149), .QN() );
  DFF_X1 cell_868_s_reg_1_s_current_state_reg ( .D(signal_1304), .CK(
        signal_1676), .Q(signal_1206), .QN() );
  DFF_X1 cell_870_s_reg_0_s_current_state_reg ( .D(signal_1054), .CK(
        signal_1676), .Q(signal_1150), .QN() );
  DFF_X1 cell_870_s_reg_1_s_current_state_reg ( .D(signal_1301), .CK(
        signal_1676), .Q(signal_1203), .QN() );
  DFF_X1 cell_872_s_reg_0_s_current_state_reg ( .D(signal_1055), .CK(
        signal_1676), .Q(signal_1151), .QN() );
  DFF_X1 cell_872_s_reg_1_s_current_state_reg ( .D(signal_1298), .CK(
        signal_1676), .Q(signal_1200), .QN() );
  DFF_X1 cell_874_s_reg_0_s_current_state_reg ( .D(signal_1056), .CK(
        signal_1676), .Q(signal_1152), .QN() );
  DFF_X1 cell_874_s_reg_1_s_current_state_reg ( .D(signal_1295), .CK(
        signal_1676), .Q(signal_1197), .QN() );
  DFF_X1 cell_876_s_reg_0_s_current_state_reg ( .D(signal_1057), .CK(
        signal_1676), .Q(signal_1153), .QN() );
  DFF_X1 cell_876_s_reg_1_s_current_state_reg ( .D(signal_1292), .CK(
        signal_1676), .Q(signal_1194), .QN() );
  DFF_X1 cell_878_s_reg_0_s_current_state_reg ( .D(signal_1058), .CK(
        signal_1676), .Q(signal_1154), .QN() );
  DFF_X1 cell_878_s_reg_1_s_current_state_reg ( .D(signal_1289), .CK(
        signal_1676), .Q(signal_1191), .QN() );
  DFF_X1 cell_880_s_reg_0_s_current_state_reg ( .D(signal_1059), .CK(
        signal_1676), .Q(signal_1155), .QN() );
  DFF_X1 cell_880_s_reg_1_s_current_state_reg ( .D(signal_1286), .CK(
        signal_1676), .Q(signal_1188), .QN() );
  DFF_X1 cell_882_s_reg_0_s_current_state_reg ( .D(signal_1060), .CK(
        signal_1676), .Q(signal_1156), .QN() );
  DFF_X1 cell_882_s_reg_1_s_current_state_reg ( .D(signal_1283), .CK(
        signal_1676), .Q(signal_1185), .QN() );
  DFF_X1 cell_884_s_reg_0_s_current_state_reg ( .D(signal_1061), .CK(
        signal_1676), .Q(signal_1157), .QN() );
  DFF_X1 cell_884_s_reg_1_s_current_state_reg ( .D(signal_1280), .CK(
        signal_1676), .Q(signal_1182), .QN() );
  DFF_X1 cell_886_s_reg_0_s_current_state_reg ( .D(signal_1062), .CK(
        signal_1676), .Q(signal_1158), .QN() );
  DFF_X1 cell_886_s_reg_1_s_current_state_reg ( .D(signal_1277), .CK(
        signal_1676), .Q(signal_1179), .QN() );
  DFF_X1 cell_888_s_reg_0_s_current_state_reg ( .D(signal_1063), .CK(
        signal_1676), .Q(signal_1159), .QN() );
  DFF_X1 cell_888_s_reg_1_s_current_state_reg ( .D(signal_1274), .CK(
        signal_1676), .Q(signal_1176), .QN() );
  DFF_X1 cell_890_s_reg_0_s_current_state_reg ( .D(signal_1064), .CK(
        signal_1676), .Q(signal_1160), .QN() );
  DFF_X1 cell_890_s_reg_1_s_current_state_reg ( .D(signal_1271), .CK(
        signal_1676), .Q(signal_1173), .QN() );
  DFF_X1 cell_892_s_reg_0_s_current_state_reg ( .D(signal_1065), .CK(
        signal_1676), .Q(signal_1161), .QN() );
  DFF_X1 cell_892_s_reg_1_s_current_state_reg ( .D(signal_1268), .CK(
        signal_1676), .Q(signal_1170), .QN() );
  DFF_X1 cell_894_s_reg_0_s_current_state_reg ( .D(signal_1066), .CK(
        signal_1676), .Q(signal_1162), .QN() );
  DFF_X1 cell_894_s_reg_1_s_current_state_reg ( .D(signal_1265), .CK(
        signal_1676), .Q(signal_1167), .QN() );
  DFF_X1 cell_896_s_reg_0_s_current_state_reg ( .D(signal_1067), .CK(
        signal_1676), .Q(signal_1163), .QN() );
  DFF_X1 cell_896_s_reg_1_s_current_state_reg ( .D(signal_1262), .CK(
        signal_1676), .Q(signal_1164), .QN() );
  DFF_X1 cell_898_s_reg_0_s_current_state_reg ( .D(signal_1068), .CK(
        signal_1676), .Q(signal_1108), .QN() );
  DFF_X1 cell_898_s_reg_1_s_current_state_reg ( .D(signal_1259), .CK(
        signal_1676), .Q(signal_1329), .QN() );
  DFF_X1 cell_900_s_reg_0_s_current_state_reg ( .D(signal_1069), .CK(
        signal_1676), .Q(signal_1109), .QN() );
  DFF_X1 cell_900_s_reg_1_s_current_state_reg ( .D(signal_1256), .CK(
        signal_1676), .Q(signal_1326), .QN() );
  DFF_X1 cell_902_s_reg_0_s_current_state_reg ( .D(signal_1070), .CK(
        signal_1676), .Q(signal_1110), .QN() );
  DFF_X1 cell_902_s_reg_1_s_current_state_reg ( .D(signal_1253), .CK(
        signal_1676), .Q(signal_1323), .QN() );
  DFF_X1 cell_904_s_reg_0_s_current_state_reg ( .D(signal_1071), .CK(
        signal_1676), .Q(signal_1111), .QN() );
  DFF_X1 cell_904_s_reg_1_s_current_state_reg ( .D(signal_1250), .CK(
        signal_1676), .Q(signal_1320), .QN() );
  DFF_X1 cell_906_s_reg_0_s_current_state_reg ( .D(signal_1072), .CK(
        signal_1676), .Q(signal_1100), .QN() );
  DFF_X1 cell_906_s_reg_1_s_current_state_reg ( .D(signal_1247), .CK(
        signal_1676), .Q(signal_1353), .QN() );
  DFF_X1 cell_908_s_reg_0_s_current_state_reg ( .D(signal_1073), .CK(
        signal_1676), .Q(signal_1101), .QN() );
  DFF_X1 cell_908_s_reg_1_s_current_state_reg ( .D(signal_1244), .CK(
        signal_1676), .Q(signal_1350), .QN() );
  DFF_X1 cell_910_s_reg_0_s_current_state_reg ( .D(signal_1074), .CK(
        signal_1676), .Q(signal_1102), .QN() );
  DFF_X1 cell_910_s_reg_1_s_current_state_reg ( .D(signal_1241), .CK(
        signal_1676), .Q(signal_1347), .QN() );
  DFF_X1 cell_912_s_reg_0_s_current_state_reg ( .D(signal_1075), .CK(
        signal_1676), .Q(signal_1103), .QN() );
  DFF_X1 cell_912_s_reg_1_s_current_state_reg ( .D(signal_1238), .CK(
        signal_1676), .Q(signal_1344), .QN() );
  DFF_X1 cell_914_s_reg_0_s_current_state_reg ( .D(signal_1076), .CK(
        signal_1676), .Q(signal_1116), .QN() );
  DFF_X1 cell_914_s_reg_1_s_current_state_reg ( .D(signal_1235), .CK(
        signal_1676), .Q(signal_1305), .QN() );
  DFF_X1 cell_916_s_reg_0_s_current_state_reg ( .D(signal_1077), .CK(
        signal_1676), .Q(signal_1117), .QN() );
  DFF_X1 cell_916_s_reg_1_s_current_state_reg ( .D(signal_1232), .CK(
        signal_1676), .Q(signal_1302), .QN() );
  DFF_X1 cell_918_s_reg_0_s_current_state_reg ( .D(signal_1078), .CK(
        signal_1676), .Q(signal_1118), .QN() );
  DFF_X1 cell_918_s_reg_1_s_current_state_reg ( .D(signal_1229), .CK(
        signal_1676), .Q(signal_1299), .QN() );
  DFF_X1 cell_920_s_reg_0_s_current_state_reg ( .D(signal_1079), .CK(
        signal_1676), .Q(signal_1119), .QN() );
  DFF_X1 cell_920_s_reg_1_s_current_state_reg ( .D(signal_1226), .CK(
        signal_1676), .Q(signal_1296), .QN() );
  DFF_X1 cell_922_s_reg_0_s_current_state_reg ( .D(signal_1080), .CK(
        signal_1676), .Q(signal_1128), .QN() );
  DFF_X1 cell_922_s_reg_1_s_current_state_reg ( .D(signal_1223), .CK(
        signal_1676), .Q(signal_1269), .QN() );
  DFF_X1 cell_924_s_reg_0_s_current_state_reg ( .D(signal_1081), .CK(
        signal_1676), .Q(signal_1129), .QN() );
  DFF_X1 cell_924_s_reg_1_s_current_state_reg ( .D(signal_1220), .CK(
        signal_1676), .Q(signal_1266), .QN() );
  DFF_X1 cell_926_s_reg_0_s_current_state_reg ( .D(signal_1082), .CK(
        signal_1676), .Q(signal_1130), .QN() );
  DFF_X1 cell_926_s_reg_1_s_current_state_reg ( .D(signal_1217), .CK(
        signal_1676), .Q(signal_1263), .QN() );
  DFF_X1 cell_928_s_reg_0_s_current_state_reg ( .D(signal_1083), .CK(
        signal_1676), .Q(signal_1131), .QN() );
  DFF_X1 cell_928_s_reg_1_s_current_state_reg ( .D(signal_1214), .CK(
        signal_1676), .Q(signal_1260), .QN() );
  DFF_X1 cell_930_s_reg_0_s_current_state_reg ( .D(signal_1084), .CK(
        signal_1676), .Q(signal_1124), .QN() );
  DFF_X1 cell_930_s_reg_1_s_current_state_reg ( .D(signal_1211), .CK(
        signal_1676), .Q(signal_1281), .QN() );
  DFF_X1 cell_932_s_reg_0_s_current_state_reg ( .D(signal_1085), .CK(
        signal_1676), .Q(signal_1125), .QN() );
  DFF_X1 cell_932_s_reg_1_s_current_state_reg ( .D(signal_1208), .CK(
        signal_1676), .Q(signal_1278), .QN() );
  DFF_X1 cell_934_s_reg_0_s_current_state_reg ( .D(signal_1086), .CK(
        signal_1676), .Q(signal_1126), .QN() );
  DFF_X1 cell_934_s_reg_1_s_current_state_reg ( .D(signal_1205), .CK(
        signal_1676), .Q(signal_1275), .QN() );
  DFF_X1 cell_936_s_reg_0_s_current_state_reg ( .D(signal_1087), .CK(
        signal_1676), .Q(signal_1127), .QN() );
  DFF_X1 cell_936_s_reg_1_s_current_state_reg ( .D(signal_1202), .CK(
        signal_1676), .Q(signal_1272), .QN() );
  DFF_X1 cell_938_s_reg_0_s_current_state_reg ( .D(signal_1088), .CK(
        signal_1676), .Q(signal_1112), .QN() );
  DFF_X1 cell_938_s_reg_1_s_current_state_reg ( .D(signal_1199), .CK(
        signal_1676), .Q(signal_1317), .QN() );
  DFF_X1 cell_940_s_reg_0_s_current_state_reg ( .D(signal_1089), .CK(
        signal_1676), .Q(signal_1113), .QN() );
  DFF_X1 cell_940_s_reg_1_s_current_state_reg ( .D(signal_1196), .CK(
        signal_1676), .Q(signal_1314), .QN() );
  DFF_X1 cell_942_s_reg_0_s_current_state_reg ( .D(signal_1090), .CK(
        signal_1676), .Q(signal_1114), .QN() );
  DFF_X1 cell_942_s_reg_1_s_current_state_reg ( .D(signal_1193), .CK(
        signal_1676), .Q(signal_1311), .QN() );
  DFF_X1 cell_944_s_reg_0_s_current_state_reg ( .D(signal_1091), .CK(
        signal_1676), .Q(signal_1115), .QN() );
  DFF_X1 cell_944_s_reg_1_s_current_state_reg ( .D(signal_1190), .CK(
        signal_1676), .Q(signal_1308), .QN() );
  DFF_X1 cell_946_s_reg_0_s_current_state_reg ( .D(signal_1092), .CK(
        signal_1676), .Q(signal_1120), .QN() );
  DFF_X1 cell_946_s_reg_1_s_current_state_reg ( .D(signal_1187), .CK(
        signal_1676), .Q(signal_1293), .QN() );
  DFF_X1 cell_948_s_reg_0_s_current_state_reg ( .D(signal_1093), .CK(
        signal_1676), .Q(signal_1121), .QN() );
  DFF_X1 cell_948_s_reg_1_s_current_state_reg ( .D(signal_1184), .CK(
        signal_1676), .Q(signal_1290), .QN() );
  DFF_X1 cell_950_s_reg_0_s_current_state_reg ( .D(signal_1094), .CK(
        signal_1676), .Q(signal_1122), .QN() );
  DFF_X1 cell_950_s_reg_1_s_current_state_reg ( .D(signal_1181), .CK(
        signal_1676), .Q(signal_1287), .QN() );
  DFF_X1 cell_952_s_reg_0_s_current_state_reg ( .D(signal_1095), .CK(
        signal_1676), .Q(signal_1123), .QN() );
  DFF_X1 cell_952_s_reg_1_s_current_state_reg ( .D(signal_1178), .CK(
        signal_1676), .Q(signal_1284), .QN() );
  DFF_X1 cell_954_s_reg_0_s_current_state_reg ( .D(signal_1096), .CK(
        signal_1676), .Q(signal_1104), .QN() );
  DFF_X1 cell_954_s_reg_1_s_current_state_reg ( .D(signal_1175), .CK(
        signal_1676), .Q(signal_1341), .QN() );
  DFF_X1 cell_956_s_reg_0_s_current_state_reg ( .D(signal_1097), .CK(
        signal_1676), .Q(signal_1105), .QN() );
  DFF_X1 cell_956_s_reg_1_s_current_state_reg ( .D(signal_1172), .CK(
        signal_1676), .Q(signal_1338), .QN() );
  DFF_X1 cell_958_s_reg_0_s_current_state_reg ( .D(signal_1098), .CK(
        signal_1676), .Q(signal_1106), .QN() );
  DFF_X1 cell_958_s_reg_1_s_current_state_reg ( .D(signal_1169), .CK(
        signal_1676), .Q(signal_1335), .QN() );
  DFF_X1 cell_960_s_reg_0_s_current_state_reg ( .D(signal_1099), .CK(
        signal_1676), .Q(signal_1107), .QN() );
  DFF_X1 cell_960_s_reg_1_s_current_state_reg ( .D(signal_1166), .CK(
        signal_1676), .Q(signal_1332), .QN() );
endmodule

