/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module Midori64_GHPC_ANF_Pipeline_d1 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, DataIn_s1, Fresh, DataOut_s0, done, DataOut_s1);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [63:0] DataIn_s1 ;
    input [63:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1458 ;
    wire signal_1461 ;
    wire signal_1464 ;
    wire signal_1467 ;
    wire signal_1470 ;
    wire signal_1473 ;
    wire signal_1476 ;
    wire signal_1479 ;
    wire signal_1482 ;
    wire signal_1485 ;
    wire signal_1488 ;
    wire signal_1491 ;
    wire signal_1494 ;
    wire signal_1497 ;
    wire signal_1500 ;
    wire signal_1503 ;
    wire signal_1506 ;
    wire signal_1509 ;
    wire signal_1512 ;
    wire signal_1515 ;
    wire signal_1518 ;
    wire signal_1521 ;
    wire signal_1524 ;
    wire signal_1527 ;
    wire signal_1530 ;
    wire signal_1533 ;
    wire signal_1536 ;
    wire signal_1539 ;
    wire signal_1542 ;
    wire signal_1545 ;
    wire signal_1548 ;
    wire signal_1551 ;
    wire signal_1554 ;
    wire signal_1557 ;
    wire signal_1560 ;
    wire signal_1563 ;
    wire signal_1566 ;
    wire signal_1569 ;
    wire signal_1572 ;
    wire signal_1575 ;
    wire signal_1578 ;
    wire signal_1581 ;
    wire signal_1584 ;
    wire signal_1587 ;
    wire signal_1590 ;
    wire signal_1593 ;
    wire signal_1596 ;
    wire signal_1599 ;
    wire signal_1602 ;
    wire signal_1605 ;
    wire signal_1608 ;
    wire signal_1611 ;
    wire signal_1614 ;
    wire signal_1617 ;
    wire signal_1620 ;
    wire signal_1623 ;
    wire signal_1626 ;
    wire signal_1629 ;
    wire signal_1632 ;
    wire signal_1635 ;
    wire signal_1638 ;
    wire signal_1641 ;
    wire signal_1644 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1662 ;
    wire signal_1664 ;
    wire signal_1666 ;
    wire signal_1668 ;
    wire signal_1670 ;
    wire signal_1672 ;
    wire signal_1674 ;
    wire signal_1676 ;
    wire signal_1678 ;
    wire signal_1680 ;
    wire signal_1682 ;
    wire signal_1684 ;
    wire signal_1686 ;
    wire signal_1688 ;
    wire signal_1690 ;
    wire signal_1692 ;
    wire signal_1694 ;
    wire signal_1696 ;
    wire signal_1698 ;
    wire signal_1700 ;
    wire signal_1702 ;
    wire signal_1704 ;
    wire signal_1706 ;
    wire signal_1708 ;
    wire signal_1710 ;
    wire signal_1712 ;
    wire signal_1714 ;
    wire signal_1716 ;
    wire signal_1718 ;
    wire signal_1720 ;
    wire signal_1722 ;
    wire signal_1724 ;
    wire signal_1726 ;
    wire signal_1728 ;
    wire signal_1730 ;
    wire signal_1732 ;
    wire signal_1734 ;
    wire signal_1736 ;
    wire signal_1738 ;
    wire signal_1740 ;
    wire signal_1742 ;
    wire signal_1744 ;
    wire signal_1746 ;
    wire signal_1748 ;
    wire signal_1750 ;
    wire signal_1752 ;
    wire signal_1754 ;
    wire signal_1756 ;
    wire signal_1758 ;
    wire signal_1760 ;
    wire signal_1762 ;
    wire signal_1764 ;
    wire signal_1766 ;
    wire signal_1768 ;
    wire signal_1770 ;
    wire signal_1772 ;
    wire signal_1774 ;
    wire signal_1776 ;
    wire signal_1778 ;
    wire signal_1780 ;
    wire signal_1782 ;
    wire signal_1784 ;
    wire signal_1786 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2528 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;

    /* cells in depth 0 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_0 ( .a ({key_s1[73], key_s0[73]}), .b ({key_s1[9], key_s0[9]}), .c ({signal_1458, signal_914}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1 ( .a ({key_s1[72], key_s0[72]}), .b ({key_s1[8], key_s0[8]}), .c ({signal_1461, signal_915}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2 ( .a ({key_s1[71], key_s0[71]}), .b ({key_s1[7], key_s0[7]}), .c ({signal_1464, signal_916}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3 ( .a ({key_s1[6], key_s0[6]}), .b ({key_s1[70], key_s0[70]}), .c ({signal_1467, signal_917}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_4 ( .a ({key_s1[127], key_s0[127]}), .b ({key_s1[63], key_s0[63]}), .c ({signal_1470, signal_860}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_5 ( .a ({key_s1[126], key_s0[126]}), .b ({key_s1[62], key_s0[62]}), .c ({signal_1473, signal_861}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_6 ( .a ({key_s1[125], key_s0[125]}), .b ({key_s1[61], key_s0[61]}), .c ({signal_1476, signal_862}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_7 ( .a ({key_s1[124], key_s0[124]}), .b ({key_s1[60], key_s0[60]}), .c ({signal_1479, signal_863}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_8 ( .a ({key_s1[5], key_s0[5]}), .b ({key_s1[69], key_s0[69]}), .c ({signal_1482, signal_918}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_9 ( .a ({key_s1[123], key_s0[123]}), .b ({key_s1[59], key_s0[59]}), .c ({signal_1485, signal_864}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_10 ( .a ({key_s1[122], key_s0[122]}), .b ({key_s1[58], key_s0[58]}), .c ({signal_1488, signal_865}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_11 ( .a ({key_s1[121], key_s0[121]}), .b ({key_s1[57], key_s0[57]}), .c ({signal_1491, signal_866}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_12 ( .a ({key_s1[120], key_s0[120]}), .b ({key_s1[56], key_s0[56]}), .c ({signal_1494, signal_867}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_13 ( .a ({key_s1[119], key_s0[119]}), .b ({key_s1[55], key_s0[55]}), .c ({signal_1497, signal_868}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_14 ( .a ({key_s1[118], key_s0[118]}), .b ({key_s1[54], key_s0[54]}), .c ({signal_1500, signal_869}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_15 ( .a ({key_s1[117], key_s0[117]}), .b ({key_s1[53], key_s0[53]}), .c ({signal_1503, signal_870}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_16 ( .a ({key_s1[116], key_s0[116]}), .b ({key_s1[52], key_s0[52]}), .c ({signal_1506, signal_871}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_17 ( .a ({key_s1[115], key_s0[115]}), .b ({key_s1[51], key_s0[51]}), .c ({signal_1509, signal_872}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_18 ( .a ({key_s1[114], key_s0[114]}), .b ({key_s1[50], key_s0[50]}), .c ({signal_1512, signal_873}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_19 ( .a ({key_s1[4], key_s0[4]}), .b ({key_s1[68], key_s0[68]}), .c ({signal_1515, signal_919}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_20 ( .a ({key_s1[113], key_s0[113]}), .b ({key_s1[49], key_s0[49]}), .c ({signal_1518, signal_874}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_21 ( .a ({key_s1[112], key_s0[112]}), .b ({key_s1[48], key_s0[48]}), .c ({signal_1521, signal_875}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_22 ( .a ({key_s1[111], key_s0[111]}), .b ({key_s1[47], key_s0[47]}), .c ({signal_1524, signal_876}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_23 ( .a ({key_s1[110], key_s0[110]}), .b ({key_s1[46], key_s0[46]}), .c ({signal_1527, signal_877}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_24 ( .a ({key_s1[109], key_s0[109]}), .b ({key_s1[45], key_s0[45]}), .c ({signal_1530, signal_878}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_25 ( .a ({key_s1[108], key_s0[108]}), .b ({key_s1[44], key_s0[44]}), .c ({signal_1533, signal_879}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_26 ( .a ({key_s1[107], key_s0[107]}), .b ({key_s1[43], key_s0[43]}), .c ({signal_1536, signal_880}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_27 ( .a ({key_s1[106], key_s0[106]}), .b ({key_s1[42], key_s0[42]}), .c ({signal_1539, signal_881}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_28 ( .a ({key_s1[105], key_s0[105]}), .b ({key_s1[41], key_s0[41]}), .c ({signal_1542, signal_882}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_29 ( .a ({key_s1[104], key_s0[104]}), .b ({key_s1[40], key_s0[40]}), .c ({signal_1545, signal_883}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_30 ( .a ({key_s1[3], key_s0[3]}), .b ({key_s1[67], key_s0[67]}), .c ({signal_1548, signal_920}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_31 ( .a ({key_s1[103], key_s0[103]}), .b ({key_s1[39], key_s0[39]}), .c ({signal_1551, signal_884}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_32 ( .a ({key_s1[102], key_s0[102]}), .b ({key_s1[38], key_s0[38]}), .c ({signal_1554, signal_885}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_33 ( .a ({key_s1[101], key_s0[101]}), .b ({key_s1[37], key_s0[37]}), .c ({signal_1557, signal_886}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_34 ( .a ({key_s1[100], key_s0[100]}), .b ({key_s1[36], key_s0[36]}), .c ({signal_1560, signal_887}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_35 ( .a ({key_s1[35], key_s0[35]}), .b ({key_s1[99], key_s0[99]}), .c ({signal_1563, signal_888}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_36 ( .a ({key_s1[34], key_s0[34]}), .b ({key_s1[98], key_s0[98]}), .c ({signal_1566, signal_889}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_37 ( .a ({key_s1[33], key_s0[33]}), .b ({key_s1[97], key_s0[97]}), .c ({signal_1569, signal_890}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_38 ( .a ({key_s1[32], key_s0[32]}), .b ({key_s1[96], key_s0[96]}), .c ({signal_1572, signal_891}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_39 ( .a ({key_s1[31], key_s0[31]}), .b ({key_s1[95], key_s0[95]}), .c ({signal_1575, signal_892}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_40 ( .a ({key_s1[30], key_s0[30]}), .b ({key_s1[94], key_s0[94]}), .c ({signal_1578, signal_893}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_41 ( .a ({key_s1[2], key_s0[2]}), .b ({key_s1[66], key_s0[66]}), .c ({signal_1581, signal_921}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_42 ( .a ({key_s1[29], key_s0[29]}), .b ({key_s1[93], key_s0[93]}), .c ({signal_1584, signal_894}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_43 ( .a ({key_s1[28], key_s0[28]}), .b ({key_s1[92], key_s0[92]}), .c ({signal_1587, signal_895}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_44 ( .a ({key_s1[27], key_s0[27]}), .b ({key_s1[91], key_s0[91]}), .c ({signal_1590, signal_896}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_45 ( .a ({key_s1[26], key_s0[26]}), .b ({key_s1[90], key_s0[90]}), .c ({signal_1593, signal_897}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_46 ( .a ({key_s1[25], key_s0[25]}), .b ({key_s1[89], key_s0[89]}), .c ({signal_1596, signal_898}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_47 ( .a ({key_s1[24], key_s0[24]}), .b ({key_s1[88], key_s0[88]}), .c ({signal_1599, signal_899}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_48 ( .a ({key_s1[23], key_s0[23]}), .b ({key_s1[87], key_s0[87]}), .c ({signal_1602, signal_900}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_49 ( .a ({key_s1[22], key_s0[22]}), .b ({key_s1[86], key_s0[86]}), .c ({signal_1605, signal_901}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_50 ( .a ({key_s1[21], key_s0[21]}), .b ({key_s1[85], key_s0[85]}), .c ({signal_1608, signal_902}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_51 ( .a ({key_s1[20], key_s0[20]}), .b ({key_s1[84], key_s0[84]}), .c ({signal_1611, signal_903}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_52 ( .a ({key_s1[1], key_s0[1]}), .b ({key_s1[65], key_s0[65]}), .c ({signal_1614, signal_922}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_53 ( .a ({key_s1[19], key_s0[19]}), .b ({key_s1[83], key_s0[83]}), .c ({signal_1617, signal_904}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_54 ( .a ({key_s1[18], key_s0[18]}), .b ({key_s1[82], key_s0[82]}), .c ({signal_1620, signal_905}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_55 ( .a ({key_s1[17], key_s0[17]}), .b ({key_s1[81], key_s0[81]}), .c ({signal_1623, signal_906}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_56 ( .a ({key_s1[16], key_s0[16]}), .b ({key_s1[80], key_s0[80]}), .c ({signal_1626, signal_907}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_57 ( .a ({key_s1[15], key_s0[15]}), .b ({key_s1[79], key_s0[79]}), .c ({signal_1629, signal_908}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_58 ( .a ({key_s1[14], key_s0[14]}), .b ({key_s1[78], key_s0[78]}), .c ({signal_1632, signal_909}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_59 ( .a ({key_s1[13], key_s0[13]}), .b ({key_s1[77], key_s0[77]}), .c ({signal_1635, signal_910}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_60 ( .a ({key_s1[12], key_s0[12]}), .b ({key_s1[76], key_s0[76]}), .c ({signal_1638, signal_911}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_61 ( .a ({key_s1[11], key_s0[11]}), .b ({key_s1[75], key_s0[75]}), .c ({signal_1641, signal_912}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_62 ( .a ({key_s1[10], key_s0[10]}), .b ({key_s1[74], key_s0[74]}), .c ({signal_1644, signal_913}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_63 ( .a ({key_s1[0], key_s0[0]}), .b ({key_s1[64], key_s0[64]}), .c ({signal_1647, signal_923}) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_266), .A2 (signal_267), .ZN (signal_265) ) ;
    NAND2_X1 cell_65 ( .A1 (signal_927), .A2 (signal_926), .ZN (signal_267) ) ;
    NAND2_X1 cell_66 ( .A1 (signal_925), .A2 (signal_924), .ZN (signal_266) ) ;
    INV_X1 cell_67 ( .A (signal_268), .ZN (signal_278) ) ;
    MUX2_X1 cell_68 ( .S (signal_281), .A (signal_269), .B (signal_270), .Z (signal_268) ) ;
    NOR2_X1 cell_69 ( .A1 (reset), .A2 (signal_271), .ZN (signal_282) ) ;
    XNOR2_X1 cell_70 ( .A (signal_927), .B (signal_926), .ZN (signal_271) ) ;
    MUX2_X1 cell_71 ( .S (signal_924), .A (signal_272), .B (signal_273), .Z (signal_280) ) ;
    NAND2_X1 cell_72 ( .A1 (signal_269), .A2 (signal_274), .ZN (signal_273) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_281), .A2 (signal_277), .ZN (signal_274) ) ;
    NOR2_X1 cell_74 ( .A1 (signal_275), .A2 (signal_283), .ZN (signal_269) ) ;
    NOR2_X1 cell_75 ( .A1 (signal_926), .A2 (reset), .ZN (signal_275) ) ;
    NOR2_X1 cell_76 ( .A1 (signal_281), .A2 (signal_270), .ZN (signal_272) ) ;
    NAND2_X1 cell_77 ( .A1 (signal_926), .A2 (signal_276), .ZN (signal_270) ) ;
    NOR2_X1 cell_78 ( .A1 (reset), .A2 (signal_279), .ZN (signal_276) ) ;
    NOR2_X1 cell_79 ( .A1 (reset), .A2 (signal_927), .ZN (signal_283) ) ;
    INV_X1 cell_80 ( .A (reset), .ZN (signal_277) ) ;
    INV_X1 cell_81 ( .A (signal_927), .ZN (signal_279) ) ;
    INV_X1 cell_85 ( .A (signal_925), .ZN (signal_281) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_153 ( .a ({signal_1458, signal_914}), .b ({DataIn_s1[9], DataIn_s0[9]}), .c ({signal_1662, signal_982}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_154 ( .a ({signal_1461, signal_915}), .b ({DataIn_s1[8], DataIn_s0[8]}), .c ({signal_1664, signal_983}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_155 ( .a ({signal_1464, signal_916}), .b ({DataIn_s1[7], DataIn_s0[7]}), .c ({signal_1666, signal_984}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_156 ( .a ({signal_1467, signal_917}), .b ({DataIn_s1[6], DataIn_s0[6]}), .c ({signal_1668, signal_985}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_157 ( .a ({signal_1470, signal_860}), .b ({DataIn_s1[63], DataIn_s0[63]}), .c ({signal_1670, signal_928}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_158 ( .a ({signal_1473, signal_861}), .b ({DataIn_s1[62], DataIn_s0[62]}), .c ({signal_1672, signal_929}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_159 ( .a ({signal_1476, signal_862}), .b ({DataIn_s1[61], DataIn_s0[61]}), .c ({signal_1674, signal_930}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_160 ( .a ({signal_1479, signal_863}), .b ({DataIn_s1[60], DataIn_s0[60]}), .c ({signal_1676, signal_931}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_161 ( .a ({signal_1482, signal_918}), .b ({DataIn_s1[5], DataIn_s0[5]}), .c ({signal_1678, signal_986}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_162 ( .a ({signal_1485, signal_864}), .b ({DataIn_s1[59], DataIn_s0[59]}), .c ({signal_1680, signal_932}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_163 ( .a ({signal_1488, signal_865}), .b ({DataIn_s1[58], DataIn_s0[58]}), .c ({signal_1682, signal_933}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_164 ( .a ({signal_1491, signal_866}), .b ({DataIn_s1[57], DataIn_s0[57]}), .c ({signal_1684, signal_934}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_165 ( .a ({signal_1494, signal_867}), .b ({DataIn_s1[56], DataIn_s0[56]}), .c ({signal_1686, signal_935}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_166 ( .a ({signal_1497, signal_868}), .b ({DataIn_s1[55], DataIn_s0[55]}), .c ({signal_1688, signal_936}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_167 ( .a ({signal_1500, signal_869}), .b ({DataIn_s1[54], DataIn_s0[54]}), .c ({signal_1690, signal_937}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_168 ( .a ({signal_1503, signal_870}), .b ({DataIn_s1[53], DataIn_s0[53]}), .c ({signal_1692, signal_938}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_169 ( .a ({signal_1506, signal_871}), .b ({DataIn_s1[52], DataIn_s0[52]}), .c ({signal_1694, signal_939}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_170 ( .a ({signal_1509, signal_872}), .b ({DataIn_s1[51], DataIn_s0[51]}), .c ({signal_1696, signal_940}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_171 ( .a ({signal_1512, signal_873}), .b ({DataIn_s1[50], DataIn_s0[50]}), .c ({signal_1698, signal_941}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_172 ( .a ({signal_1515, signal_919}), .b ({DataIn_s1[4], DataIn_s0[4]}), .c ({signal_1700, signal_987}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_173 ( .a ({signal_1518, signal_874}), .b ({DataIn_s1[49], DataIn_s0[49]}), .c ({signal_1702, signal_942}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_174 ( .a ({signal_1521, signal_875}), .b ({DataIn_s1[48], DataIn_s0[48]}), .c ({signal_1704, signal_943}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_175 ( .a ({signal_1524, signal_876}), .b ({DataIn_s1[47], DataIn_s0[47]}), .c ({signal_1706, signal_944}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_176 ( .a ({signal_1527, signal_877}), .b ({DataIn_s1[46], DataIn_s0[46]}), .c ({signal_1708, signal_945}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_177 ( .a ({signal_1530, signal_878}), .b ({DataIn_s1[45], DataIn_s0[45]}), .c ({signal_1710, signal_946}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_178 ( .a ({signal_1533, signal_879}), .b ({DataIn_s1[44], DataIn_s0[44]}), .c ({signal_1712, signal_947}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_179 ( .a ({signal_1536, signal_880}), .b ({DataIn_s1[43], DataIn_s0[43]}), .c ({signal_1714, signal_948}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_180 ( .a ({signal_1539, signal_881}), .b ({DataIn_s1[42], DataIn_s0[42]}), .c ({signal_1716, signal_949}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_181 ( .a ({signal_1542, signal_882}), .b ({DataIn_s1[41], DataIn_s0[41]}), .c ({signal_1718, signal_950}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_182 ( .a ({signal_1545, signal_883}), .b ({DataIn_s1[40], DataIn_s0[40]}), .c ({signal_1720, signal_951}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_183 ( .a ({signal_1548, signal_920}), .b ({DataIn_s1[3], DataIn_s0[3]}), .c ({signal_1722, signal_988}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_184 ( .a ({signal_1551, signal_884}), .b ({DataIn_s1[39], DataIn_s0[39]}), .c ({signal_1724, signal_952}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_185 ( .a ({signal_1554, signal_885}), .b ({DataIn_s1[38], DataIn_s0[38]}), .c ({signal_1726, signal_953}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_186 ( .a ({signal_1557, signal_886}), .b ({DataIn_s1[37], DataIn_s0[37]}), .c ({signal_1728, signal_954}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_187 ( .a ({signal_1560, signal_887}), .b ({DataIn_s1[36], DataIn_s0[36]}), .c ({signal_1730, signal_955}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_188 ( .a ({signal_1563, signal_888}), .b ({DataIn_s1[35], DataIn_s0[35]}), .c ({signal_1732, signal_956}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_189 ( .a ({signal_1566, signal_889}), .b ({DataIn_s1[34], DataIn_s0[34]}), .c ({signal_1734, signal_957}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_190 ( .a ({signal_1569, signal_890}), .b ({DataIn_s1[33], DataIn_s0[33]}), .c ({signal_1736, signal_958}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_191 ( .a ({signal_1572, signal_891}), .b ({DataIn_s1[32], DataIn_s0[32]}), .c ({signal_1738, signal_959}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_192 ( .a ({signal_1575, signal_892}), .b ({DataIn_s1[31], DataIn_s0[31]}), .c ({signal_1740, signal_960}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_193 ( .a ({signal_1578, signal_893}), .b ({DataIn_s1[30], DataIn_s0[30]}), .c ({signal_1742, signal_961}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_194 ( .a ({signal_1581, signal_921}), .b ({DataIn_s1[2], DataIn_s0[2]}), .c ({signal_1744, signal_989}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_195 ( .a ({signal_1584, signal_894}), .b ({DataIn_s1[29], DataIn_s0[29]}), .c ({signal_1746, signal_962}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_196 ( .a ({signal_1587, signal_895}), .b ({DataIn_s1[28], DataIn_s0[28]}), .c ({signal_1748, signal_963}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_197 ( .a ({signal_1590, signal_896}), .b ({DataIn_s1[27], DataIn_s0[27]}), .c ({signal_1750, signal_964}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_198 ( .a ({signal_1593, signal_897}), .b ({DataIn_s1[26], DataIn_s0[26]}), .c ({signal_1752, signal_965}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_199 ( .a ({signal_1596, signal_898}), .b ({DataIn_s1[25], DataIn_s0[25]}), .c ({signal_1754, signal_966}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_200 ( .a ({signal_1599, signal_899}), .b ({DataIn_s1[24], DataIn_s0[24]}), .c ({signal_1756, signal_967}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_201 ( .a ({signal_1602, signal_900}), .b ({DataIn_s1[23], DataIn_s0[23]}), .c ({signal_1758, signal_968}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_202 ( .a ({signal_1605, signal_901}), .b ({DataIn_s1[22], DataIn_s0[22]}), .c ({signal_1760, signal_969}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_203 ( .a ({signal_1608, signal_902}), .b ({DataIn_s1[21], DataIn_s0[21]}), .c ({signal_1762, signal_970}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_204 ( .a ({signal_1611, signal_903}), .b ({DataIn_s1[20], DataIn_s0[20]}), .c ({signal_1764, signal_971}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_205 ( .a ({signal_1614, signal_922}), .b ({DataIn_s1[1], DataIn_s0[1]}), .c ({signal_1766, signal_990}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_206 ( .a ({signal_1617, signal_904}), .b ({DataIn_s1[19], DataIn_s0[19]}), .c ({signal_1768, signal_972}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_207 ( .a ({signal_1620, signal_905}), .b ({DataIn_s1[18], DataIn_s0[18]}), .c ({signal_1770, signal_973}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_208 ( .a ({signal_1623, signal_906}), .b ({DataIn_s1[17], DataIn_s0[17]}), .c ({signal_1772, signal_974}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_209 ( .a ({signal_1626, signal_907}), .b ({DataIn_s1[16], DataIn_s0[16]}), .c ({signal_1774, signal_975}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_210 ( .a ({signal_1629, signal_908}), .b ({DataIn_s1[15], DataIn_s0[15]}), .c ({signal_1776, signal_976}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_211 ( .a ({signal_1632, signal_909}), .b ({DataIn_s1[14], DataIn_s0[14]}), .c ({signal_1778, signal_977}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_212 ( .a ({signal_1635, signal_910}), .b ({DataIn_s1[13], DataIn_s0[13]}), .c ({signal_1780, signal_978}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_213 ( .a ({signal_1638, signal_911}), .b ({DataIn_s1[12], DataIn_s0[12]}), .c ({signal_1782, signal_979}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_214 ( .a ({signal_1641, signal_912}), .b ({DataIn_s1[11], DataIn_s0[11]}), .c ({signal_1784, signal_980}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_215 ( .a ({signal_1644, signal_913}), .b ({DataIn_s1[10], DataIn_s0[10]}), .c ({signal_1786, signal_981}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_216 ( .a ({signal_1647, signal_923}), .b ({DataIn_s1[0], DataIn_s0[0]}), .c ({signal_1788, signal_991}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_283 ( .a ({signal_1653, signal_310}), .b ({1'b0, signal_1453}), .c ({signal_2254, signal_286}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_290 ( .a ({signal_2038, signal_362}), .b ({1'b0, signal_1440}), .c ({signal_2310, signal_287}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_296 ( .a ({signal_2034, signal_358}), .b ({1'b0, signal_1441}), .c ({signal_2311, signal_288}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_301 ( .a ({signal_2030, signal_354}), .b ({1'b0, signal_1442}), .c ({signal_2312, signal_289}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_305 ( .a ({signal_1652, signal_306}), .b ({1'b0, signal_1454}), .c ({signal_2313, signal_290}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_308 ( .a ({signal_2026, signal_350}), .b ({1'b0, signal_1443}), .c ({signal_2378, signal_291}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_313 ( .a ({signal_2022, signal_346}), .b ({1'b0, signal_1444}), .c ({signal_2255, signal_292}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_318 ( .a ({signal_2018, signal_342}), .b ({1'b0, signal_1445}), .c ({signal_2314, signal_293}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_324 ( .a ({signal_2014, signal_338}), .b ({1'b0, signal_1446}), .c ({signal_2256, signal_294}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_329 ( .a ({signal_2010, signal_334}), .b ({1'b0, signal_1447}), .c ({signal_2315, signal_295}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_335 ( .a ({signal_2006, signal_330}), .b ({1'b0, signal_1448}), .c ({signal_2372, signal_296}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_340 ( .a ({signal_2003, signal_326}), .b ({1'b0, signal_1449}), .c ({signal_2316, signal_297}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_345 ( .a ({signal_1999, signal_322}), .b ({1'b0, signal_1450}), .c ({signal_2257, signal_298}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_351 ( .a ({signal_1995, signal_318}), .b ({1'b0, signal_1451}), .c ({signal_2317, signal_299}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_356 ( .a ({signal_1994, signal_314}), .b ({1'b0, signal_1452}), .c ({signal_2318, signal_300}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_360 ( .a ({signal_1648, signal_302}), .b ({1'b0, signal_1455}), .c ({signal_2319, signal_301}) ) ;
    NAND2_X1 cell_361 ( .A1 (signal_366), .A2 (signal_367), .ZN (signal_1446) ) ;
    NOR2_X1 cell_362 ( .A1 (signal_368), .A2 (signal_369), .ZN (signal_366) ) ;
    OR2_X1 cell_363 ( .A1 (signal_370), .A2 (signal_371), .ZN (signal_369) ) ;
    NAND2_X1 cell_364 ( .A1 (signal_372), .A2 (signal_373), .ZN (signal_1447) ) ;
    NAND2_X1 cell_365 ( .A1 (signal_374), .A2 (signal_375), .ZN (signal_1448) ) ;
    NOR2_X1 cell_366 ( .A1 (signal_1444), .A2 (signal_376), .ZN (signal_375) ) ;
    NAND2_X1 cell_367 ( .A1 (signal_377), .A2 (signal_378), .ZN (signal_376) ) ;
    NOR2_X1 cell_368 ( .A1 (signal_379), .A2 (signal_380), .ZN (signal_377) ) ;
    NAND2_X1 cell_369 ( .A1 (signal_381), .A2 (signal_382), .ZN (signal_1449) ) ;
    NOR2_X1 cell_370 ( .A1 (signal_383), .A2 (signal_384), .ZN (signal_382) ) ;
    NAND2_X1 cell_371 ( .A1 (signal_385), .A2 (signal_386), .ZN (signal_1450) ) ;
    NOR2_X1 cell_372 ( .A1 (signal_371), .A2 (signal_387), .ZN (signal_386) ) ;
    NAND2_X1 cell_373 ( .A1 (signal_388), .A2 (signal_378), .ZN (signal_387) ) ;
    NAND2_X1 cell_374 ( .A1 (signal_389), .A2 (signal_388), .ZN (signal_1451) ) ;
    NOR2_X1 cell_375 ( .A1 (signal_390), .A2 (signal_391), .ZN (signal_388) ) ;
    NAND2_X1 cell_376 ( .A1 (signal_392), .A2 (signal_393), .ZN (signal_1452) ) ;
    NOR2_X1 cell_377 ( .A1 (signal_368), .A2 (signal_394), .ZN (signal_392) ) ;
    NAND2_X1 cell_378 ( .A1 (signal_395), .A2 (signal_378), .ZN (signal_394) ) ;
    INV_X1 cell_379 ( .A (signal_396), .ZN (signal_395) ) ;
    OR2_X1 cell_380 ( .A1 (signal_368), .A2 (signal_397), .ZN (signal_1453) ) ;
    NAND2_X1 cell_381 ( .A1 (signal_381), .A2 (signal_398), .ZN (signal_397) ) ;
    NOR2_X1 cell_382 ( .A1 (signal_399), .A2 (signal_371), .ZN (signal_381) ) ;
    NAND2_X1 cell_383 ( .A1 (signal_400), .A2 (signal_373), .ZN (signal_368) ) ;
    NAND2_X1 cell_384 ( .A1 (signal_401), .A2 (signal_402), .ZN (signal_1454) ) ;
    NOR2_X1 cell_385 ( .A1 (signal_396), .A2 (signal_403), .ZN (signal_402) ) ;
    OR2_X1 cell_386 ( .A1 (signal_371), .A2 (signal_379), .ZN (signal_403) ) ;
    INV_X1 cell_387 ( .A (signal_400), .ZN (signal_379) ) ;
    NAND2_X1 cell_388 ( .A1 (signal_404), .A2 (signal_405), .ZN (signal_400) ) ;
    NAND2_X1 cell_389 ( .A1 (signal_406), .A2 (signal_407), .ZN (signal_405) ) ;
    NOR2_X1 cell_390 ( .A1 (signal_455), .A2 (signal_408), .ZN (signal_371) ) ;
    MUX2_X1 cell_391 ( .S (signal_925), .A (signal_409), .B (signal_410), .Z (signal_408) ) ;
    NAND2_X1 cell_392 ( .A1 (signal_411), .A2 (signal_412), .ZN (signal_1440) ) ;
    NOR2_X1 cell_393 ( .A1 (signal_383), .A2 (signal_396), .ZN (signal_411) ) ;
    NAND2_X1 cell_394 ( .A1 (signal_413), .A2 (signal_389), .ZN (signal_1441) ) ;
    NOR2_X1 cell_395 ( .A1 (signal_414), .A2 (signal_415), .ZN (signal_389) ) ;
    NAND2_X1 cell_396 ( .A1 (signal_367), .A2 (signal_378), .ZN (signal_415) ) ;
    OR2_X1 cell_397 ( .A1 (signal_454), .A2 (signal_416), .ZN (signal_378) ) ;
    MUX2_X1 cell_398 ( .S (signal_925), .A (signal_417), .B (signal_418), .Z (signal_416) ) ;
    NAND2_X1 cell_399 ( .A1 (signal_398), .A2 (signal_419), .ZN (signal_1442) ) ;
    NOR2_X1 cell_400 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_419) ) ;
    INV_X1 cell_401 ( .A (signal_413), .ZN (signal_421) ) ;
    NOR2_X1 cell_402 ( .A1 (signal_422), .A2 (signal_391), .ZN (signal_398) ) ;
    NAND2_X1 cell_403 ( .A1 (signal_423), .A2 (signal_393), .ZN (signal_1443) ) ;
    INV_X1 cell_404 ( .A (signal_399), .ZN (signal_393) ) ;
    NOR2_X1 cell_405 ( .A1 (signal_380), .A2 (signal_424), .ZN (signal_423) ) ;
    NAND2_X1 cell_406 ( .A1 (signal_372), .A2 (signal_413), .ZN (signal_424) ) ;
    NOR2_X1 cell_407 ( .A1 (signal_390), .A2 (signal_414), .ZN (signal_372) ) ;
    NAND2_X1 cell_408 ( .A1 (signal_385), .A2 (signal_425), .ZN (signal_414) ) ;
    NAND2_X1 cell_409 ( .A1 (signal_454), .A2 (signal_426), .ZN (signal_425) ) ;
    NAND2_X1 cell_410 ( .A1 (signal_418), .A2 (signal_406), .ZN (signal_426) ) ;
    NOR2_X1 cell_411 ( .A1 (signal_383), .A2 (signal_427), .ZN (signal_385) ) ;
    NOR2_X1 cell_412 ( .A1 (signal_455), .A2 (signal_428), .ZN (signal_427) ) ;
    MUX2_X1 cell_413 ( .S (signal_925), .A (signal_407), .B (signal_417), .Z (signal_428) ) ;
    NOR2_X1 cell_414 ( .A1 (signal_454), .A2 (signal_429), .ZN (signal_383) ) ;
    MUX2_X1 cell_415 ( .S (signal_925), .A (signal_409), .B (signal_430), .Z (signal_429) ) ;
    OR2_X1 cell_416 ( .A1 (signal_384), .A2 (signal_370), .ZN (signal_1444) ) ;
    NAND2_X1 cell_417 ( .A1 (signal_413), .A2 (signal_373), .ZN (signal_384) ) ;
    NAND2_X1 cell_418 ( .A1 (signal_431), .A2 (signal_432), .ZN (signal_373) ) ;
    AND2_X1 cell_419 ( .A1 (signal_455), .A2 (signal_925), .ZN (signal_432) ) ;
    NOR2_X1 cell_420 ( .A1 (signal_433), .A2 (signal_396), .ZN (signal_413) ) ;
    NOR2_X1 cell_421 ( .A1 (signal_454), .A2 (signal_434), .ZN (signal_396) ) ;
    MUX2_X1 cell_422 ( .S (signal_925), .A (signal_418), .B (signal_417), .Z (signal_434) ) ;
    NOR2_X1 cell_423 ( .A1 (signal_454), .A2 (signal_435), .ZN (signal_433) ) ;
    MUX2_X1 cell_424 ( .S (signal_925), .A (signal_430), .B (signal_409), .Z (signal_435) ) ;
    NAND2_X1 cell_425 ( .A1 (signal_436), .A2 (signal_412), .ZN (signal_1445) ) ;
    NOR2_X1 cell_426 ( .A1 (signal_437), .A2 (signal_370), .ZN (signal_412) ) ;
    NOR2_X1 cell_427 ( .A1 (signal_455), .A2 (signal_438), .ZN (signal_370) ) ;
    MUX2_X1 cell_428 ( .S (signal_925), .A (signal_418), .B (signal_406), .Z (signal_438) ) ;
    INV_X1 cell_429 ( .A (signal_439), .ZN (signal_437) ) ;
    INV_X1 cell_430 ( .A (signal_390), .ZN (signal_436) ) ;
    NAND2_X1 cell_431 ( .A1 (signal_401), .A2 (signal_439), .ZN (signal_1455) ) ;
    NOR2_X1 cell_432 ( .A1 (signal_380), .A2 (signal_391), .ZN (signal_439) ) ;
    NOR2_X1 cell_433 ( .A1 (signal_455), .A2 (signal_440), .ZN (signal_391) ) ;
    MUX2_X1 cell_434 ( .S (signal_925), .A (signal_410), .B (signal_409), .Z (signal_440) ) ;
    NAND2_X1 cell_435 ( .A1 (signal_441), .A2 (signal_442), .ZN (signal_409) ) ;
    NAND2_X1 cell_436 ( .A1 (signal_443), .A2 (signal_926), .ZN (signal_410) ) ;
    NOR2_X1 cell_437 ( .A1 (signal_455), .A2 (signal_444), .ZN (signal_380) ) ;
    MUX2_X1 cell_438 ( .S (signal_925), .A (signal_417), .B (signal_407), .Z (signal_444) ) ;
    NAND2_X1 cell_439 ( .A1 (enc_dec), .A2 (signal_431), .ZN (signal_407) ) ;
    NOR2_X1 cell_440 ( .A1 (signal_924), .A2 (signal_442), .ZN (signal_431) ) ;
    NAND2_X1 cell_441 ( .A1 (signal_445), .A2 (signal_442), .ZN (signal_417) ) ;
    NOR2_X1 cell_442 ( .A1 (signal_399), .A2 (signal_446), .ZN (signal_401) ) ;
    NAND2_X1 cell_443 ( .A1 (signal_374), .A2 (signal_367), .ZN (signal_446) ) ;
    NAND2_X1 cell_444 ( .A1 (signal_420), .A2 (signal_447), .ZN (signal_367) ) ;
    OR2_X1 cell_445 ( .A1 (signal_443), .A2 (signal_441), .ZN (signal_447) ) ;
    AND2_X1 cell_446 ( .A1 (signal_926), .A2 (signal_404), .ZN (signal_420) ) ;
    NOR2_X1 cell_447 ( .A1 (signal_454), .A2 (signal_925), .ZN (signal_404) ) ;
    NOR2_X1 cell_448 ( .A1 (signal_390), .A2 (signal_422), .ZN (signal_374) ) ;
    NOR2_X1 cell_449 ( .A1 (signal_455), .A2 (signal_448), .ZN (signal_422) ) ;
    MUX2_X1 cell_450 ( .S (signal_925), .A (signal_406), .B (signal_418), .Z (signal_448) ) ;
    NAND2_X1 cell_451 ( .A1 (enc_dec), .A2 (signal_449), .ZN (signal_418) ) ;
    NOR2_X1 cell_452 ( .A1 (signal_924), .A2 (signal_926), .ZN (signal_449) ) ;
    NAND2_X1 cell_453 ( .A1 (signal_926), .A2 (signal_445), .ZN (signal_406) ) ;
    NOR2_X1 cell_454 ( .A1 (enc_dec), .A2 (signal_450), .ZN (signal_445) ) ;
    INV_X1 cell_455 ( .A (signal_924), .ZN (signal_450) ) ;
    NOR2_X1 cell_456 ( .A1 (signal_455), .A2 (signal_451), .ZN (signal_390) ) ;
    MUX2_X1 cell_457 ( .S (signal_925), .A (signal_430), .B (signal_452), .Z (signal_451) ) ;
    NOR2_X1 cell_458 ( .A1 (signal_455), .A2 (signal_453), .ZN (signal_399) ) ;
    MUX2_X1 cell_459 ( .S (signal_925), .A (signal_452), .B (signal_430), .Z (signal_453) ) ;
    NAND2_X1 cell_460 ( .A1 (signal_443), .A2 (signal_442), .ZN (signal_430) ) ;
    INV_X1 cell_461 ( .A (signal_926), .ZN (signal_442) ) ;
    NOR2_X1 cell_462 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_443) ) ;
    NAND2_X1 cell_463 ( .A1 (signal_441), .A2 (signal_926), .ZN (signal_452) ) ;
    AND2_X1 cell_464 ( .A1 (enc_dec), .A2 (signal_924), .ZN (signal_441) ) ;
    INV_X1 cell_465 ( .A (signal_454), .ZN (signal_455) ) ;
    INV_X1 cell_466 ( .A (signal_927), .ZN (signal_454) ) ;
    INV_X1 cell_467 ( .A (signal_927), .ZN (signal_456) ) ;
    INV_X1 cell_468 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_469 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_470 ( .A (signal_456), .ZN (signal_457) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_471 ( .s (signal_927), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1648, signal_302}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_472 ( .s (signal_927), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1649, signal_303}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_473 ( .s (signal_927), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1650, signal_304}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_474 ( .s (signal_927), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1651, signal_305}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_475 ( .s (signal_927), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1652, signal_306}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_476 ( .s (signal_459), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1991, signal_307}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_477 ( .s (signal_457), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1992, signal_308}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_478 ( .s (signal_458), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1993, signal_309}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_479 ( .s (signal_927), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1653, signal_310}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_480 ( .s (signal_927), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1654, signal_311}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_481 ( .s (signal_927), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1655, signal_312}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_482 ( .s (signal_927), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1656, signal_313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_483 ( .s (signal_458), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1994, signal_314}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_484 ( .s (signal_927), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1657, signal_315}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_485 ( .s (signal_927), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1658, signal_316}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_486 ( .s (signal_927), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1659, signal_317}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_487 ( .s (signal_457), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1995, signal_318}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_488 ( .s (signal_459), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1996, signal_319}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_489 ( .s (signal_457), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1997, signal_320}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_490 ( .s (signal_457), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1998, signal_321}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_491 ( .s (signal_457), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1999, signal_322}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_492 ( .s (signal_457), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_2000, signal_323}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_493 ( .s (signal_458), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_2001, signal_324}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_494 ( .s (signal_459), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_2002, signal_325}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_495 ( .s (signal_457), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_2003, signal_326}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_496 ( .s (signal_458), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_2004, signal_327}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_497 ( .s (signal_927), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1660, signal_328}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_498 ( .s (signal_457), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_2005, signal_329}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_499 ( .s (signal_457), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_2006, signal_330}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_500 ( .s (signal_457), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_2007, signal_331}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_501 ( .s (signal_457), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_2008, signal_332}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_502 ( .s (signal_457), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_2009, signal_333}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_503 ( .s (signal_457), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_2010, signal_334}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_504 ( .s (signal_457), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_2011, signal_335}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_505 ( .s (signal_457), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_2012, signal_336}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_506 ( .s (signal_457), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_2013, signal_337}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_507 ( .s (signal_457), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_2014, signal_338}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_508 ( .s (signal_457), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_2015, signal_339}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_509 ( .s (signal_457), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_2016, signal_340}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_510 ( .s (signal_457), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_2017, signal_341}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_511 ( .s (signal_458), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_2018, signal_342}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_512 ( .s (signal_458), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_2019, signal_343}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_513 ( .s (signal_458), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_2020, signal_344}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_514 ( .s (signal_458), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_2021, signal_345}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_515 ( .s (signal_458), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_2022, signal_346}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_516 ( .s (signal_458), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_2023, signal_347}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_517 ( .s (signal_458), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_2024, signal_348}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_518 ( .s (signal_458), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_2025, signal_349}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_519 ( .s (signal_458), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_2026, signal_350}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_520 ( .s (signal_458), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_2027, signal_351}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_521 ( .s (signal_458), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_2028, signal_352}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_522 ( .s (signal_458), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_2029, signal_353}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_523 ( .s (signal_459), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_2030, signal_354}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_524 ( .s (signal_459), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_2031, signal_355}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_525 ( .s (signal_459), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_2032, signal_356}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_526 ( .s (signal_459), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_2033, signal_357}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_527 ( .s (signal_459), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_2034, signal_358}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_528 ( .s (signal_459), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_2035, signal_359}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_529 ( .s (signal_459), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_2036, signal_360}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_530 ( .s (signal_459), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_2037, signal_361}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_531 ( .s (signal_459), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_2038, signal_362}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_532 ( .s (signal_459), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_2039, signal_363}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_533 ( .s (signal_459), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_2040, signal_364}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_534 ( .s (signal_459), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_2041, signal_365}) ) ;

    /* cells in depth 1 */
    buf_clk cell_1256 ( .C (clk), .D (signal_265), .Q (signal_2528) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_914), .Q (signal_2530) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_1458), .Q (signal_2532) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_915), .Q (signal_2534) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_1461), .Q (signal_2536) ) ;
    buf_clk cell_1266 ( .C (clk), .D (signal_916), .Q (signal_2538) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_1464), .Q (signal_2540) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_917), .Q (signal_2542) ) ;
    buf_clk cell_1272 ( .C (clk), .D (signal_1467), .Q (signal_2544) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_860), .Q (signal_2546) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_1470), .Q (signal_2548) ) ;
    buf_clk cell_1278 ( .C (clk), .D (signal_861), .Q (signal_2550) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_1473), .Q (signal_2552) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_862), .Q (signal_2554) ) ;
    buf_clk cell_1284 ( .C (clk), .D (signal_1476), .Q (signal_2556) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_863), .Q (signal_2558) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_1479), .Q (signal_2560) ) ;
    buf_clk cell_1290 ( .C (clk), .D (signal_918), .Q (signal_2562) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_1482), .Q (signal_2564) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_864), .Q (signal_2566) ) ;
    buf_clk cell_1296 ( .C (clk), .D (signal_1485), .Q (signal_2568) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_865), .Q (signal_2570) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_1488), .Q (signal_2572) ) ;
    buf_clk cell_1302 ( .C (clk), .D (signal_866), .Q (signal_2574) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_1491), .Q (signal_2576) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_867), .Q (signal_2578) ) ;
    buf_clk cell_1308 ( .C (clk), .D (signal_1494), .Q (signal_2580) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_868), .Q (signal_2582) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_1497), .Q (signal_2584) ) ;
    buf_clk cell_1314 ( .C (clk), .D (signal_869), .Q (signal_2586) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_1500), .Q (signal_2588) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_870), .Q (signal_2590) ) ;
    buf_clk cell_1320 ( .C (clk), .D (signal_1503), .Q (signal_2592) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_871), .Q (signal_2594) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_1506), .Q (signal_2596) ) ;
    buf_clk cell_1326 ( .C (clk), .D (signal_872), .Q (signal_2598) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_1509), .Q (signal_2600) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_873), .Q (signal_2602) ) ;
    buf_clk cell_1332 ( .C (clk), .D (signal_1512), .Q (signal_2604) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_919), .Q (signal_2606) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_1515), .Q (signal_2608) ) ;
    buf_clk cell_1338 ( .C (clk), .D (signal_874), .Q (signal_2610) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_1518), .Q (signal_2612) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_875), .Q (signal_2614) ) ;
    buf_clk cell_1344 ( .C (clk), .D (signal_1521), .Q (signal_2616) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_876), .Q (signal_2618) ) ;
    buf_clk cell_1348 ( .C (clk), .D (signal_1524), .Q (signal_2620) ) ;
    buf_clk cell_1350 ( .C (clk), .D (signal_877), .Q (signal_2622) ) ;
    buf_clk cell_1352 ( .C (clk), .D (signal_1527), .Q (signal_2624) ) ;
    buf_clk cell_1354 ( .C (clk), .D (signal_878), .Q (signal_2626) ) ;
    buf_clk cell_1356 ( .C (clk), .D (signal_1530), .Q (signal_2628) ) ;
    buf_clk cell_1358 ( .C (clk), .D (signal_879), .Q (signal_2630) ) ;
    buf_clk cell_1360 ( .C (clk), .D (signal_1533), .Q (signal_2632) ) ;
    buf_clk cell_1362 ( .C (clk), .D (signal_880), .Q (signal_2634) ) ;
    buf_clk cell_1364 ( .C (clk), .D (signal_1536), .Q (signal_2636) ) ;
    buf_clk cell_1366 ( .C (clk), .D (signal_881), .Q (signal_2638) ) ;
    buf_clk cell_1368 ( .C (clk), .D (signal_1539), .Q (signal_2640) ) ;
    buf_clk cell_1370 ( .C (clk), .D (signal_882), .Q (signal_2642) ) ;
    buf_clk cell_1372 ( .C (clk), .D (signal_1542), .Q (signal_2644) ) ;
    buf_clk cell_1374 ( .C (clk), .D (signal_883), .Q (signal_2646) ) ;
    buf_clk cell_1376 ( .C (clk), .D (signal_1545), .Q (signal_2648) ) ;
    buf_clk cell_1378 ( .C (clk), .D (signal_920), .Q (signal_2650) ) ;
    buf_clk cell_1380 ( .C (clk), .D (signal_1548), .Q (signal_2652) ) ;
    buf_clk cell_1382 ( .C (clk), .D (signal_884), .Q (signal_2654) ) ;
    buf_clk cell_1384 ( .C (clk), .D (signal_1551), .Q (signal_2656) ) ;
    buf_clk cell_1386 ( .C (clk), .D (signal_885), .Q (signal_2658) ) ;
    buf_clk cell_1388 ( .C (clk), .D (signal_1554), .Q (signal_2660) ) ;
    buf_clk cell_1390 ( .C (clk), .D (signal_886), .Q (signal_2662) ) ;
    buf_clk cell_1392 ( .C (clk), .D (signal_1557), .Q (signal_2664) ) ;
    buf_clk cell_1394 ( .C (clk), .D (signal_887), .Q (signal_2666) ) ;
    buf_clk cell_1396 ( .C (clk), .D (signal_1560), .Q (signal_2668) ) ;
    buf_clk cell_1398 ( .C (clk), .D (signal_888), .Q (signal_2670) ) ;
    buf_clk cell_1400 ( .C (clk), .D (signal_1563), .Q (signal_2672) ) ;
    buf_clk cell_1402 ( .C (clk), .D (signal_889), .Q (signal_2674) ) ;
    buf_clk cell_1404 ( .C (clk), .D (signal_1566), .Q (signal_2676) ) ;
    buf_clk cell_1406 ( .C (clk), .D (signal_890), .Q (signal_2678) ) ;
    buf_clk cell_1408 ( .C (clk), .D (signal_1569), .Q (signal_2680) ) ;
    buf_clk cell_1410 ( .C (clk), .D (signal_891), .Q (signal_2682) ) ;
    buf_clk cell_1412 ( .C (clk), .D (signal_1572), .Q (signal_2684) ) ;
    buf_clk cell_1414 ( .C (clk), .D (signal_892), .Q (signal_2686) ) ;
    buf_clk cell_1416 ( .C (clk), .D (signal_1575), .Q (signal_2688) ) ;
    buf_clk cell_1418 ( .C (clk), .D (signal_893), .Q (signal_2690) ) ;
    buf_clk cell_1420 ( .C (clk), .D (signal_1578), .Q (signal_2692) ) ;
    buf_clk cell_1422 ( .C (clk), .D (signal_921), .Q (signal_2694) ) ;
    buf_clk cell_1424 ( .C (clk), .D (signal_1581), .Q (signal_2696) ) ;
    buf_clk cell_1426 ( .C (clk), .D (signal_894), .Q (signal_2698) ) ;
    buf_clk cell_1428 ( .C (clk), .D (signal_1584), .Q (signal_2700) ) ;
    buf_clk cell_1430 ( .C (clk), .D (signal_895), .Q (signal_2702) ) ;
    buf_clk cell_1432 ( .C (clk), .D (signal_1587), .Q (signal_2704) ) ;
    buf_clk cell_1434 ( .C (clk), .D (signal_896), .Q (signal_2706) ) ;
    buf_clk cell_1436 ( .C (clk), .D (signal_1590), .Q (signal_2708) ) ;
    buf_clk cell_1438 ( .C (clk), .D (signal_897), .Q (signal_2710) ) ;
    buf_clk cell_1440 ( .C (clk), .D (signal_1593), .Q (signal_2712) ) ;
    buf_clk cell_1442 ( .C (clk), .D (signal_898), .Q (signal_2714) ) ;
    buf_clk cell_1444 ( .C (clk), .D (signal_1596), .Q (signal_2716) ) ;
    buf_clk cell_1446 ( .C (clk), .D (signal_899), .Q (signal_2718) ) ;
    buf_clk cell_1448 ( .C (clk), .D (signal_1599), .Q (signal_2720) ) ;
    buf_clk cell_1450 ( .C (clk), .D (signal_900), .Q (signal_2722) ) ;
    buf_clk cell_1452 ( .C (clk), .D (signal_1602), .Q (signal_2724) ) ;
    buf_clk cell_1454 ( .C (clk), .D (signal_901), .Q (signal_2726) ) ;
    buf_clk cell_1456 ( .C (clk), .D (signal_1605), .Q (signal_2728) ) ;
    buf_clk cell_1458 ( .C (clk), .D (signal_902), .Q (signal_2730) ) ;
    buf_clk cell_1460 ( .C (clk), .D (signal_1608), .Q (signal_2732) ) ;
    buf_clk cell_1462 ( .C (clk), .D (signal_903), .Q (signal_2734) ) ;
    buf_clk cell_1464 ( .C (clk), .D (signal_1611), .Q (signal_2736) ) ;
    buf_clk cell_1466 ( .C (clk), .D (signal_922), .Q (signal_2738) ) ;
    buf_clk cell_1468 ( .C (clk), .D (signal_1614), .Q (signal_2740) ) ;
    buf_clk cell_1470 ( .C (clk), .D (signal_904), .Q (signal_2742) ) ;
    buf_clk cell_1472 ( .C (clk), .D (signal_1617), .Q (signal_2744) ) ;
    buf_clk cell_1474 ( .C (clk), .D (signal_905), .Q (signal_2746) ) ;
    buf_clk cell_1476 ( .C (clk), .D (signal_1620), .Q (signal_2748) ) ;
    buf_clk cell_1478 ( .C (clk), .D (signal_906), .Q (signal_2750) ) ;
    buf_clk cell_1480 ( .C (clk), .D (signal_1623), .Q (signal_2752) ) ;
    buf_clk cell_1482 ( .C (clk), .D (signal_907), .Q (signal_2754) ) ;
    buf_clk cell_1484 ( .C (clk), .D (signal_1626), .Q (signal_2756) ) ;
    buf_clk cell_1486 ( .C (clk), .D (signal_908), .Q (signal_2758) ) ;
    buf_clk cell_1488 ( .C (clk), .D (signal_1629), .Q (signal_2760) ) ;
    buf_clk cell_1490 ( .C (clk), .D (signal_909), .Q (signal_2762) ) ;
    buf_clk cell_1492 ( .C (clk), .D (signal_1632), .Q (signal_2764) ) ;
    buf_clk cell_1494 ( .C (clk), .D (signal_910), .Q (signal_2766) ) ;
    buf_clk cell_1496 ( .C (clk), .D (signal_1635), .Q (signal_2768) ) ;
    buf_clk cell_1498 ( .C (clk), .D (signal_911), .Q (signal_2770) ) ;
    buf_clk cell_1500 ( .C (clk), .D (signal_1638), .Q (signal_2772) ) ;
    buf_clk cell_1502 ( .C (clk), .D (signal_912), .Q (signal_2774) ) ;
    buf_clk cell_1504 ( .C (clk), .D (signal_1641), .Q (signal_2776) ) ;
    buf_clk cell_1506 ( .C (clk), .D (signal_913), .Q (signal_2778) ) ;
    buf_clk cell_1508 ( .C (clk), .D (signal_1644), .Q (signal_2780) ) ;
    buf_clk cell_1510 ( .C (clk), .D (signal_923), .Q (signal_2782) ) ;
    buf_clk cell_1512 ( .C (clk), .D (signal_1647), .Q (signal_2784) ) ;
    buf_clk cell_1514 ( .C (clk), .D (signal_311), .Q (signal_2786) ) ;
    buf_clk cell_1516 ( .C (clk), .D (signal_1654), .Q (signal_2788) ) ;
    buf_clk cell_1518 ( .C (clk), .D (signal_286), .Q (signal_2790) ) ;
    buf_clk cell_1520 ( .C (clk), .D (signal_2254), .Q (signal_2792) ) ;
    buf_clk cell_1522 ( .C (clk), .D (signal_309), .Q (signal_2794) ) ;
    buf_clk cell_1524 ( .C (clk), .D (signal_1993), .Q (signal_2796) ) ;
    buf_clk cell_1526 ( .C (clk), .D (signal_308), .Q (signal_2798) ) ;
    buf_clk cell_1528 ( .C (clk), .D (signal_1992), .Q (signal_2800) ) ;
    buf_clk cell_1530 ( .C (clk), .D (signal_365), .Q (signal_2802) ) ;
    buf_clk cell_1532 ( .C (clk), .D (signal_2041), .Q (signal_2804) ) ;
    buf_clk cell_1534 ( .C (clk), .D (signal_364), .Q (signal_2806) ) ;
    buf_clk cell_1536 ( .C (clk), .D (signal_2040), .Q (signal_2808) ) ;
    buf_clk cell_1538 ( .C (clk), .D (signal_363), .Q (signal_2810) ) ;
    buf_clk cell_1540 ( .C (clk), .D (signal_2039), .Q (signal_2812) ) ;
    buf_clk cell_1542 ( .C (clk), .D (signal_287), .Q (signal_2814) ) ;
    buf_clk cell_1544 ( .C (clk), .D (signal_2310), .Q (signal_2816) ) ;
    buf_clk cell_1546 ( .C (clk), .D (signal_307), .Q (signal_2818) ) ;
    buf_clk cell_1548 ( .C (clk), .D (signal_1991), .Q (signal_2820) ) ;
    buf_clk cell_1550 ( .C (clk), .D (signal_361), .Q (signal_2822) ) ;
    buf_clk cell_1552 ( .C (clk), .D (signal_2037), .Q (signal_2824) ) ;
    buf_clk cell_1554 ( .C (clk), .D (signal_360), .Q (signal_2826) ) ;
    buf_clk cell_1556 ( .C (clk), .D (signal_2036), .Q (signal_2828) ) ;
    buf_clk cell_1558 ( .C (clk), .D (signal_359), .Q (signal_2830) ) ;
    buf_clk cell_1560 ( .C (clk), .D (signal_2035), .Q (signal_2832) ) ;
    buf_clk cell_1562 ( .C (clk), .D (signal_288), .Q (signal_2834) ) ;
    buf_clk cell_1564 ( .C (clk), .D (signal_2311), .Q (signal_2836) ) ;
    buf_clk cell_1566 ( .C (clk), .D (signal_357), .Q (signal_2838) ) ;
    buf_clk cell_1568 ( .C (clk), .D (signal_2033), .Q (signal_2840) ) ;
    buf_clk cell_1570 ( .C (clk), .D (signal_356), .Q (signal_2842) ) ;
    buf_clk cell_1572 ( .C (clk), .D (signal_2032), .Q (signal_2844) ) ;
    buf_clk cell_1574 ( .C (clk), .D (signal_355), .Q (signal_2846) ) ;
    buf_clk cell_1576 ( .C (clk), .D (signal_2031), .Q (signal_2848) ) ;
    buf_clk cell_1578 ( .C (clk), .D (signal_289), .Q (signal_2850) ) ;
    buf_clk cell_1580 ( .C (clk), .D (signal_2312), .Q (signal_2852) ) ;
    buf_clk cell_1582 ( .C (clk), .D (signal_353), .Q (signal_2854) ) ;
    buf_clk cell_1584 ( .C (clk), .D (signal_2029), .Q (signal_2856) ) ;
    buf_clk cell_1586 ( .C (clk), .D (signal_352), .Q (signal_2858) ) ;
    buf_clk cell_1588 ( .C (clk), .D (signal_2028), .Q (signal_2860) ) ;
    buf_clk cell_1590 ( .C (clk), .D (signal_290), .Q (signal_2862) ) ;
    buf_clk cell_1592 ( .C (clk), .D (signal_2313), .Q (signal_2864) ) ;
    buf_clk cell_1594 ( .C (clk), .D (signal_351), .Q (signal_2866) ) ;
    buf_clk cell_1596 ( .C (clk), .D (signal_2027), .Q (signal_2868) ) ;
    buf_clk cell_1598 ( .C (clk), .D (signal_291), .Q (signal_2870) ) ;
    buf_clk cell_1600 ( .C (clk), .D (signal_2378), .Q (signal_2872) ) ;
    buf_clk cell_1602 ( .C (clk), .D (signal_349), .Q (signal_2874) ) ;
    buf_clk cell_1604 ( .C (clk), .D (signal_2025), .Q (signal_2876) ) ;
    buf_clk cell_1606 ( .C (clk), .D (signal_348), .Q (signal_2878) ) ;
    buf_clk cell_1608 ( .C (clk), .D (signal_2024), .Q (signal_2880) ) ;
    buf_clk cell_1610 ( .C (clk), .D (signal_347), .Q (signal_2882) ) ;
    buf_clk cell_1612 ( .C (clk), .D (signal_2023), .Q (signal_2884) ) ;
    buf_clk cell_1614 ( .C (clk), .D (signal_292), .Q (signal_2886) ) ;
    buf_clk cell_1616 ( .C (clk), .D (signal_2255), .Q (signal_2888) ) ;
    buf_clk cell_1618 ( .C (clk), .D (signal_345), .Q (signal_2890) ) ;
    buf_clk cell_1620 ( .C (clk), .D (signal_2021), .Q (signal_2892) ) ;
    buf_clk cell_1622 ( .C (clk), .D (signal_344), .Q (signal_2894) ) ;
    buf_clk cell_1624 ( .C (clk), .D (signal_2020), .Q (signal_2896) ) ;
    buf_clk cell_1626 ( .C (clk), .D (signal_343), .Q (signal_2898) ) ;
    buf_clk cell_1628 ( .C (clk), .D (signal_2019), .Q (signal_2900) ) ;
    buf_clk cell_1630 ( .C (clk), .D (signal_293), .Q (signal_2902) ) ;
    buf_clk cell_1632 ( .C (clk), .D (signal_2314), .Q (signal_2904) ) ;
    buf_clk cell_1634 ( .C (clk), .D (signal_305), .Q (signal_2906) ) ;
    buf_clk cell_1636 ( .C (clk), .D (signal_1651), .Q (signal_2908) ) ;
    buf_clk cell_1638 ( .C (clk), .D (signal_341), .Q (signal_2910) ) ;
    buf_clk cell_1640 ( .C (clk), .D (signal_2017), .Q (signal_2912) ) ;
    buf_clk cell_1642 ( .C (clk), .D (signal_340), .Q (signal_2914) ) ;
    buf_clk cell_1644 ( .C (clk), .D (signal_2016), .Q (signal_2916) ) ;
    buf_clk cell_1646 ( .C (clk), .D (signal_339), .Q (signal_2918) ) ;
    buf_clk cell_1648 ( .C (clk), .D (signal_2015), .Q (signal_2920) ) ;
    buf_clk cell_1650 ( .C (clk), .D (signal_294), .Q (signal_2922) ) ;
    buf_clk cell_1652 ( .C (clk), .D (signal_2256), .Q (signal_2924) ) ;
    buf_clk cell_1654 ( .C (clk), .D (signal_337), .Q (signal_2926) ) ;
    buf_clk cell_1656 ( .C (clk), .D (signal_2013), .Q (signal_2928) ) ;
    buf_clk cell_1658 ( .C (clk), .D (signal_336), .Q (signal_2930) ) ;
    buf_clk cell_1660 ( .C (clk), .D (signal_2012), .Q (signal_2932) ) ;
    buf_clk cell_1662 ( .C (clk), .D (signal_335), .Q (signal_2934) ) ;
    buf_clk cell_1664 ( .C (clk), .D (signal_2011), .Q (signal_2936) ) ;
    buf_clk cell_1666 ( .C (clk), .D (signal_295), .Q (signal_2938) ) ;
    buf_clk cell_1668 ( .C (clk), .D (signal_2315), .Q (signal_2940) ) ;
    buf_clk cell_1670 ( .C (clk), .D (signal_333), .Q (signal_2942) ) ;
    buf_clk cell_1672 ( .C (clk), .D (signal_2009), .Q (signal_2944) ) ;
    buf_clk cell_1674 ( .C (clk), .D (signal_332), .Q (signal_2946) ) ;
    buf_clk cell_1676 ( .C (clk), .D (signal_2008), .Q (signal_2948) ) ;
    buf_clk cell_1678 ( .C (clk), .D (signal_304), .Q (signal_2950) ) ;
    buf_clk cell_1680 ( .C (clk), .D (signal_1650), .Q (signal_2952) ) ;
    buf_clk cell_1682 ( .C (clk), .D (signal_331), .Q (signal_2954) ) ;
    buf_clk cell_1684 ( .C (clk), .D (signal_2007), .Q (signal_2956) ) ;
    buf_clk cell_1686 ( .C (clk), .D (signal_296), .Q (signal_2958) ) ;
    buf_clk cell_1688 ( .C (clk), .D (signal_2372), .Q (signal_2960) ) ;
    buf_clk cell_1690 ( .C (clk), .D (signal_329), .Q (signal_2962) ) ;
    buf_clk cell_1692 ( .C (clk), .D (signal_2005), .Q (signal_2964) ) ;
    buf_clk cell_1694 ( .C (clk), .D (signal_328), .Q (signal_2966) ) ;
    buf_clk cell_1696 ( .C (clk), .D (signal_1660), .Q (signal_2968) ) ;
    buf_clk cell_1698 ( .C (clk), .D (signal_327), .Q (signal_2970) ) ;
    buf_clk cell_1700 ( .C (clk), .D (signal_2004), .Q (signal_2972) ) ;
    buf_clk cell_1702 ( .C (clk), .D (signal_297), .Q (signal_2974) ) ;
    buf_clk cell_1704 ( .C (clk), .D (signal_2316), .Q (signal_2976) ) ;
    buf_clk cell_1706 ( .C (clk), .D (signal_325), .Q (signal_2978) ) ;
    buf_clk cell_1708 ( .C (clk), .D (signal_2002), .Q (signal_2980) ) ;
    buf_clk cell_1710 ( .C (clk), .D (signal_324), .Q (signal_2982) ) ;
    buf_clk cell_1712 ( .C (clk), .D (signal_2001), .Q (signal_2984) ) ;
    buf_clk cell_1714 ( .C (clk), .D (signal_323), .Q (signal_2986) ) ;
    buf_clk cell_1716 ( .C (clk), .D (signal_2000), .Q (signal_2988) ) ;
    buf_clk cell_1718 ( .C (clk), .D (signal_298), .Q (signal_2990) ) ;
    buf_clk cell_1720 ( .C (clk), .D (signal_2257), .Q (signal_2992) ) ;
    buf_clk cell_1722 ( .C (clk), .D (signal_303), .Q (signal_2994) ) ;
    buf_clk cell_1724 ( .C (clk), .D (signal_1649), .Q (signal_2996) ) ;
    buf_clk cell_1726 ( .C (clk), .D (signal_321), .Q (signal_2998) ) ;
    buf_clk cell_1728 ( .C (clk), .D (signal_1998), .Q (signal_3000) ) ;
    buf_clk cell_1730 ( .C (clk), .D (signal_320), .Q (signal_3002) ) ;
    buf_clk cell_1732 ( .C (clk), .D (signal_1997), .Q (signal_3004) ) ;
    buf_clk cell_1734 ( .C (clk), .D (signal_319), .Q (signal_3006) ) ;
    buf_clk cell_1736 ( .C (clk), .D (signal_1996), .Q (signal_3008) ) ;
    buf_clk cell_1738 ( .C (clk), .D (signal_299), .Q (signal_3010) ) ;
    buf_clk cell_1740 ( .C (clk), .D (signal_2317), .Q (signal_3012) ) ;
    buf_clk cell_1742 ( .C (clk), .D (signal_317), .Q (signal_3014) ) ;
    buf_clk cell_1744 ( .C (clk), .D (signal_1659), .Q (signal_3016) ) ;
    buf_clk cell_1746 ( .C (clk), .D (signal_316), .Q (signal_3018) ) ;
    buf_clk cell_1748 ( .C (clk), .D (signal_1658), .Q (signal_3020) ) ;
    buf_clk cell_1750 ( .C (clk), .D (signal_315), .Q (signal_3022) ) ;
    buf_clk cell_1752 ( .C (clk), .D (signal_1657), .Q (signal_3024) ) ;
    buf_clk cell_1754 ( .C (clk), .D (signal_300), .Q (signal_3026) ) ;
    buf_clk cell_1756 ( .C (clk), .D (signal_2318), .Q (signal_3028) ) ;
    buf_clk cell_1758 ( .C (clk), .D (signal_313), .Q (signal_3030) ) ;
    buf_clk cell_1760 ( .C (clk), .D (signal_1656), .Q (signal_3032) ) ;
    buf_clk cell_1762 ( .C (clk), .D (signal_312), .Q (signal_3034) ) ;
    buf_clk cell_1764 ( .C (clk), .D (signal_1655), .Q (signal_3036) ) ;
    buf_clk cell_1766 ( .C (clk), .D (signal_301), .Q (signal_3038) ) ;
    buf_clk cell_1768 ( .C (clk), .D (signal_2319), .Q (signal_3040) ) ;
    buf_clk cell_1770 ( .C (clk), .D (reset), .Q (signal_3042) ) ;
    buf_clk cell_1772 ( .C (clk), .D (signal_991), .Q (signal_3044) ) ;
    buf_clk cell_1774 ( .C (clk), .D (signal_1788), .Q (signal_3046) ) ;
    buf_clk cell_1776 ( .C (clk), .D (signal_990), .Q (signal_3048) ) ;
    buf_clk cell_1778 ( .C (clk), .D (signal_1766), .Q (signal_3050) ) ;
    buf_clk cell_1780 ( .C (clk), .D (signal_989), .Q (signal_3052) ) ;
    buf_clk cell_1782 ( .C (clk), .D (signal_1744), .Q (signal_3054) ) ;
    buf_clk cell_1784 ( .C (clk), .D (signal_988), .Q (signal_3056) ) ;
    buf_clk cell_1786 ( .C (clk), .D (signal_1722), .Q (signal_3058) ) ;
    buf_clk cell_1788 ( .C (clk), .D (signal_987), .Q (signal_3060) ) ;
    buf_clk cell_1790 ( .C (clk), .D (signal_1700), .Q (signal_3062) ) ;
    buf_clk cell_1792 ( .C (clk), .D (signal_986), .Q (signal_3064) ) ;
    buf_clk cell_1794 ( .C (clk), .D (signal_1678), .Q (signal_3066) ) ;
    buf_clk cell_1796 ( .C (clk), .D (signal_985), .Q (signal_3068) ) ;
    buf_clk cell_1798 ( .C (clk), .D (signal_1668), .Q (signal_3070) ) ;
    buf_clk cell_1800 ( .C (clk), .D (signal_984), .Q (signal_3072) ) ;
    buf_clk cell_1802 ( .C (clk), .D (signal_1666), .Q (signal_3074) ) ;
    buf_clk cell_1804 ( .C (clk), .D (signal_983), .Q (signal_3076) ) ;
    buf_clk cell_1806 ( .C (clk), .D (signal_1664), .Q (signal_3078) ) ;
    buf_clk cell_1808 ( .C (clk), .D (signal_982), .Q (signal_3080) ) ;
    buf_clk cell_1810 ( .C (clk), .D (signal_1662), .Q (signal_3082) ) ;
    buf_clk cell_1812 ( .C (clk), .D (signal_981), .Q (signal_3084) ) ;
    buf_clk cell_1814 ( .C (clk), .D (signal_1786), .Q (signal_3086) ) ;
    buf_clk cell_1816 ( .C (clk), .D (signal_980), .Q (signal_3088) ) ;
    buf_clk cell_1818 ( .C (clk), .D (signal_1784), .Q (signal_3090) ) ;
    buf_clk cell_1820 ( .C (clk), .D (signal_979), .Q (signal_3092) ) ;
    buf_clk cell_1822 ( .C (clk), .D (signal_1782), .Q (signal_3094) ) ;
    buf_clk cell_1824 ( .C (clk), .D (signal_978), .Q (signal_3096) ) ;
    buf_clk cell_1826 ( .C (clk), .D (signal_1780), .Q (signal_3098) ) ;
    buf_clk cell_1828 ( .C (clk), .D (signal_977), .Q (signal_3100) ) ;
    buf_clk cell_1830 ( .C (clk), .D (signal_1778), .Q (signal_3102) ) ;
    buf_clk cell_1832 ( .C (clk), .D (signal_976), .Q (signal_3104) ) ;
    buf_clk cell_1834 ( .C (clk), .D (signal_1776), .Q (signal_3106) ) ;
    buf_clk cell_1836 ( .C (clk), .D (signal_975), .Q (signal_3108) ) ;
    buf_clk cell_1838 ( .C (clk), .D (signal_1774), .Q (signal_3110) ) ;
    buf_clk cell_1840 ( .C (clk), .D (signal_974), .Q (signal_3112) ) ;
    buf_clk cell_1842 ( .C (clk), .D (signal_1772), .Q (signal_3114) ) ;
    buf_clk cell_1844 ( .C (clk), .D (signal_973), .Q (signal_3116) ) ;
    buf_clk cell_1846 ( .C (clk), .D (signal_1770), .Q (signal_3118) ) ;
    buf_clk cell_1848 ( .C (clk), .D (signal_972), .Q (signal_3120) ) ;
    buf_clk cell_1850 ( .C (clk), .D (signal_1768), .Q (signal_3122) ) ;
    buf_clk cell_1852 ( .C (clk), .D (signal_971), .Q (signal_3124) ) ;
    buf_clk cell_1854 ( .C (clk), .D (signal_1764), .Q (signal_3126) ) ;
    buf_clk cell_1856 ( .C (clk), .D (signal_970), .Q (signal_3128) ) ;
    buf_clk cell_1858 ( .C (clk), .D (signal_1762), .Q (signal_3130) ) ;
    buf_clk cell_1860 ( .C (clk), .D (signal_969), .Q (signal_3132) ) ;
    buf_clk cell_1862 ( .C (clk), .D (signal_1760), .Q (signal_3134) ) ;
    buf_clk cell_1864 ( .C (clk), .D (signal_968), .Q (signal_3136) ) ;
    buf_clk cell_1866 ( .C (clk), .D (signal_1758), .Q (signal_3138) ) ;
    buf_clk cell_1868 ( .C (clk), .D (signal_967), .Q (signal_3140) ) ;
    buf_clk cell_1870 ( .C (clk), .D (signal_1756), .Q (signal_3142) ) ;
    buf_clk cell_1872 ( .C (clk), .D (signal_966), .Q (signal_3144) ) ;
    buf_clk cell_1874 ( .C (clk), .D (signal_1754), .Q (signal_3146) ) ;
    buf_clk cell_1876 ( .C (clk), .D (signal_965), .Q (signal_3148) ) ;
    buf_clk cell_1878 ( .C (clk), .D (signal_1752), .Q (signal_3150) ) ;
    buf_clk cell_1880 ( .C (clk), .D (signal_964), .Q (signal_3152) ) ;
    buf_clk cell_1882 ( .C (clk), .D (signal_1750), .Q (signal_3154) ) ;
    buf_clk cell_1884 ( .C (clk), .D (signal_963), .Q (signal_3156) ) ;
    buf_clk cell_1886 ( .C (clk), .D (signal_1748), .Q (signal_3158) ) ;
    buf_clk cell_1888 ( .C (clk), .D (signal_962), .Q (signal_3160) ) ;
    buf_clk cell_1890 ( .C (clk), .D (signal_1746), .Q (signal_3162) ) ;
    buf_clk cell_1892 ( .C (clk), .D (signal_961), .Q (signal_3164) ) ;
    buf_clk cell_1894 ( .C (clk), .D (signal_1742), .Q (signal_3166) ) ;
    buf_clk cell_1896 ( .C (clk), .D (signal_960), .Q (signal_3168) ) ;
    buf_clk cell_1898 ( .C (clk), .D (signal_1740), .Q (signal_3170) ) ;
    buf_clk cell_1900 ( .C (clk), .D (signal_959), .Q (signal_3172) ) ;
    buf_clk cell_1902 ( .C (clk), .D (signal_1738), .Q (signal_3174) ) ;
    buf_clk cell_1904 ( .C (clk), .D (signal_958), .Q (signal_3176) ) ;
    buf_clk cell_1906 ( .C (clk), .D (signal_1736), .Q (signal_3178) ) ;
    buf_clk cell_1908 ( .C (clk), .D (signal_957), .Q (signal_3180) ) ;
    buf_clk cell_1910 ( .C (clk), .D (signal_1734), .Q (signal_3182) ) ;
    buf_clk cell_1912 ( .C (clk), .D (signal_956), .Q (signal_3184) ) ;
    buf_clk cell_1914 ( .C (clk), .D (signal_1732), .Q (signal_3186) ) ;
    buf_clk cell_1916 ( .C (clk), .D (signal_955), .Q (signal_3188) ) ;
    buf_clk cell_1918 ( .C (clk), .D (signal_1730), .Q (signal_3190) ) ;
    buf_clk cell_1920 ( .C (clk), .D (signal_954), .Q (signal_3192) ) ;
    buf_clk cell_1922 ( .C (clk), .D (signal_1728), .Q (signal_3194) ) ;
    buf_clk cell_1924 ( .C (clk), .D (signal_953), .Q (signal_3196) ) ;
    buf_clk cell_1926 ( .C (clk), .D (signal_1726), .Q (signal_3198) ) ;
    buf_clk cell_1928 ( .C (clk), .D (signal_952), .Q (signal_3200) ) ;
    buf_clk cell_1930 ( .C (clk), .D (signal_1724), .Q (signal_3202) ) ;
    buf_clk cell_1932 ( .C (clk), .D (signal_951), .Q (signal_3204) ) ;
    buf_clk cell_1934 ( .C (clk), .D (signal_1720), .Q (signal_3206) ) ;
    buf_clk cell_1936 ( .C (clk), .D (signal_950), .Q (signal_3208) ) ;
    buf_clk cell_1938 ( .C (clk), .D (signal_1718), .Q (signal_3210) ) ;
    buf_clk cell_1940 ( .C (clk), .D (signal_949), .Q (signal_3212) ) ;
    buf_clk cell_1942 ( .C (clk), .D (signal_1716), .Q (signal_3214) ) ;
    buf_clk cell_1944 ( .C (clk), .D (signal_948), .Q (signal_3216) ) ;
    buf_clk cell_1946 ( .C (clk), .D (signal_1714), .Q (signal_3218) ) ;
    buf_clk cell_1948 ( .C (clk), .D (signal_947), .Q (signal_3220) ) ;
    buf_clk cell_1950 ( .C (clk), .D (signal_1712), .Q (signal_3222) ) ;
    buf_clk cell_1952 ( .C (clk), .D (signal_946), .Q (signal_3224) ) ;
    buf_clk cell_1954 ( .C (clk), .D (signal_1710), .Q (signal_3226) ) ;
    buf_clk cell_1956 ( .C (clk), .D (signal_945), .Q (signal_3228) ) ;
    buf_clk cell_1958 ( .C (clk), .D (signal_1708), .Q (signal_3230) ) ;
    buf_clk cell_1960 ( .C (clk), .D (signal_944), .Q (signal_3232) ) ;
    buf_clk cell_1962 ( .C (clk), .D (signal_1706), .Q (signal_3234) ) ;
    buf_clk cell_1964 ( .C (clk), .D (signal_943), .Q (signal_3236) ) ;
    buf_clk cell_1966 ( .C (clk), .D (signal_1704), .Q (signal_3238) ) ;
    buf_clk cell_1968 ( .C (clk), .D (signal_942), .Q (signal_3240) ) ;
    buf_clk cell_1970 ( .C (clk), .D (signal_1702), .Q (signal_3242) ) ;
    buf_clk cell_1972 ( .C (clk), .D (signal_941), .Q (signal_3244) ) ;
    buf_clk cell_1974 ( .C (clk), .D (signal_1698), .Q (signal_3246) ) ;
    buf_clk cell_1976 ( .C (clk), .D (signal_940), .Q (signal_3248) ) ;
    buf_clk cell_1978 ( .C (clk), .D (signal_1696), .Q (signal_3250) ) ;
    buf_clk cell_1980 ( .C (clk), .D (signal_939), .Q (signal_3252) ) ;
    buf_clk cell_1982 ( .C (clk), .D (signal_1694), .Q (signal_3254) ) ;
    buf_clk cell_1984 ( .C (clk), .D (signal_938), .Q (signal_3256) ) ;
    buf_clk cell_1986 ( .C (clk), .D (signal_1692), .Q (signal_3258) ) ;
    buf_clk cell_1988 ( .C (clk), .D (signal_937), .Q (signal_3260) ) ;
    buf_clk cell_1990 ( .C (clk), .D (signal_1690), .Q (signal_3262) ) ;
    buf_clk cell_1992 ( .C (clk), .D (signal_936), .Q (signal_3264) ) ;
    buf_clk cell_1994 ( .C (clk), .D (signal_1688), .Q (signal_3266) ) ;
    buf_clk cell_1996 ( .C (clk), .D (signal_935), .Q (signal_3268) ) ;
    buf_clk cell_1998 ( .C (clk), .D (signal_1686), .Q (signal_3270) ) ;
    buf_clk cell_2000 ( .C (clk), .D (signal_934), .Q (signal_3272) ) ;
    buf_clk cell_2002 ( .C (clk), .D (signal_1684), .Q (signal_3274) ) ;
    buf_clk cell_2004 ( .C (clk), .D (signal_933), .Q (signal_3276) ) ;
    buf_clk cell_2006 ( .C (clk), .D (signal_1682), .Q (signal_3278) ) ;
    buf_clk cell_2008 ( .C (clk), .D (signal_932), .Q (signal_3280) ) ;
    buf_clk cell_2010 ( .C (clk), .D (signal_1680), .Q (signal_3282) ) ;
    buf_clk cell_2012 ( .C (clk), .D (signal_931), .Q (signal_3284) ) ;
    buf_clk cell_2014 ( .C (clk), .D (signal_1676), .Q (signal_3286) ) ;
    buf_clk cell_2016 ( .C (clk), .D (signal_930), .Q (signal_3288) ) ;
    buf_clk cell_2018 ( .C (clk), .D (signal_1674), .Q (signal_3290) ) ;
    buf_clk cell_2020 ( .C (clk), .D (signal_929), .Q (signal_3292) ) ;
    buf_clk cell_2022 ( .C (clk), .D (signal_1672), .Q (signal_3294) ) ;
    buf_clk cell_2024 ( .C (clk), .D (signal_928), .Q (signal_3296) ) ;
    buf_clk cell_2026 ( .C (clk), .D (signal_1670), .Q (signal_3298) ) ;
    buf_clk cell_2028 ( .C (clk), .D (enc_dec), .Q (signal_3300) ) ;
    buf_clk cell_2030 ( .C (clk), .D (signal_283), .Q (signal_3302) ) ;
    buf_clk cell_2032 ( .C (clk), .D (signal_282), .Q (signal_3304) ) ;
    buf_clk cell_2034 ( .C (clk), .D (signal_278), .Q (signal_3306) ) ;
    buf_clk cell_2036 ( .C (clk), .D (signal_280), .Q (signal_3308) ) ;

    /* cells in depth 2 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_89 ( .a ({signal_2533, signal_2531}), .b ({signal_1907, signal_1302}), .c ({DataOut_s1[9], DataOut_s0[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_90 ( .a ({signal_2537, signal_2535}), .b ({signal_1908, signal_1303}), .c ({DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_91 ( .a ({signal_2541, signal_2539}), .b ({signal_1869, signal_1264}), .c ({DataOut_s1[7], DataOut_s0[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_92 ( .a ({signal_2545, signal_2543}), .b ({signal_1870, signal_1265}), .c ({DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_93 ( .a ({signal_2549, signal_2547}), .b ({signal_1853, signal_1248}), .c ({DataOut_s1[63], DataOut_s0[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_94 ( .a ({signal_2553, signal_2551}), .b ({signal_1854, signal_1249}), .c ({DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_95 ( .a ({signal_2557, signal_2555}), .b ({signal_1855, signal_1250}), .c ({DataOut_s1[61], DataOut_s0[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_96 ( .a ({signal_2561, signal_2559}), .b ({signal_1856, signal_1251}), .c ({DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_97 ( .a ({signal_2565, signal_2563}), .b ({signal_1871, signal_1266}), .c ({DataOut_s1[5], DataOut_s0[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_98 ( .a ({signal_2569, signal_2567}), .b ({signal_1881, signal_1276}), .c ({DataOut_s1[59], DataOut_s0[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_99 ( .a ({signal_2573, signal_2571}), .b ({signal_1882, signal_1277}), .c ({DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_100 ( .a ({signal_2577, signal_2575}), .b ({signal_1883, signal_1278}), .c ({DataOut_s1[57], DataOut_s0[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_101 ( .a ({signal_2581, signal_2579}), .b ({signal_1884, signal_1279}), .c ({DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_102 ( .a ({signal_2585, signal_2583}), .b ({signal_1909, signal_1304}), .c ({DataOut_s1[55], DataOut_s0[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_103 ( .a ({signal_2589, signal_2587}), .b ({signal_1910, signal_1305}), .c ({DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_104 ( .a ({signal_2593, signal_2591}), .b ({signal_1911, signal_1306}), .c ({DataOut_s1[53], DataOut_s0[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_105 ( .a ({signal_2597, signal_2595}), .b ({signal_1912, signal_1307}), .c ({DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_106 ( .a ({signal_2601, signal_2599}), .b ({signal_1889, signal_1284}), .c ({DataOut_s1[51], DataOut_s0[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_107 ( .a ({signal_2605, signal_2603}), .b ({signal_1890, signal_1285}), .c ({DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_108 ( .a ({signal_2609, signal_2607}), .b ({signal_1872, signal_1267}), .c ({DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_109 ( .a ({signal_2613, signal_2611}), .b ({signal_1891, signal_1286}), .c ({DataOut_s1[49], DataOut_s0[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_110 ( .a ({signal_2617, signal_2615}), .b ({signal_1892, signal_1287}), .c ({DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_111 ( .a ({signal_2621, signal_2619}), .b ({signal_1873, signal_1268}), .c ({DataOut_s1[47], DataOut_s0[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_112 ( .a ({signal_2625, signal_2623}), .b ({signal_1874, signal_1269}), .c ({DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_113 ( .a ({signal_2629, signal_2627}), .b ({signal_1875, signal_1270}), .c ({DataOut_s1[45], DataOut_s0[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_114 ( .a ({signal_2633, signal_2631}), .b ({signal_1876, signal_1271}), .c ({DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_115 ( .a ({signal_2637, signal_2635}), .b ({signal_1861, signal_1256}), .c ({DataOut_s1[43], DataOut_s0[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_116 ( .a ({signal_2641, signal_2639}), .b ({signal_1862, signal_1257}), .c ({DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_117 ( .a ({signal_2645, signal_2643}), .b ({signal_1863, signal_1258}), .c ({DataOut_s1[41], DataOut_s0[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_118 ( .a ({signal_2649, signal_2647}), .b ({signal_1864, signal_1259}), .c ({DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_119 ( .a ({signal_2653, signal_2651}), .b ({signal_1865, signal_1260}), .c ({DataOut_s1[3], DataOut_s0[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_120 ( .a ({signal_2657, signal_2655}), .b ({signal_1897, signal_1292}), .c ({DataOut_s1[39], DataOut_s0[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_121 ( .a ({signal_2661, signal_2659}), .b ({signal_1898, signal_1293}), .c ({DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_122 ( .a ({signal_2665, signal_2663}), .b ({signal_1899, signal_1294}), .c ({DataOut_s1[37], DataOut_s0[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_123 ( .a ({signal_2669, signal_2667}), .b ({signal_1900, signal_1295}), .c ({DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_124 ( .a ({signal_2673, signal_2671}), .b ({signal_1901, signal_1296}), .c ({DataOut_s1[35], DataOut_s0[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_125 ( .a ({signal_2677, signal_2675}), .b ({signal_1902, signal_1297}), .c ({DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_126 ( .a ({signal_2681, signal_2679}), .b ({signal_1903, signal_1298}), .c ({DataOut_s1[33], DataOut_s0[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_127 ( .a ({signal_2685, signal_2683}), .b ({signal_1904, signal_1299}), .c ({DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_128 ( .a ({signal_2689, signal_2687}), .b ({signal_1913, signal_1308}), .c ({DataOut_s1[31], DataOut_s0[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_129 ( .a ({signal_2693, signal_2691}), .b ({signal_1914, signal_1309}), .c ({DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_130 ( .a ({signal_2697, signal_2695}), .b ({signal_1866, signal_1261}), .c ({DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_131 ( .a ({signal_2701, signal_2699}), .b ({signal_1915, signal_1310}), .c ({DataOut_s1[29], DataOut_s0[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_132 ( .a ({signal_2705, signal_2703}), .b ({signal_1916, signal_1311}), .c ({DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_133 ( .a ({signal_2709, signal_2707}), .b ({signal_1885, signal_1280}), .c ({DataOut_s1[27], DataOut_s0[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_134 ( .a ({signal_2713, signal_2711}), .b ({signal_1886, signal_1281}), .c ({DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_135 ( .a ({signal_2717, signal_2715}), .b ({signal_1887, signal_1282}), .c ({DataOut_s1[25], DataOut_s0[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_136 ( .a ({signal_2721, signal_2719}), .b ({signal_1888, signal_1283}), .c ({DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_137 ( .a ({signal_2725, signal_2723}), .b ({signal_1857, signal_1252}), .c ({DataOut_s1[23], DataOut_s0[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_138 ( .a ({signal_2729, signal_2727}), .b ({signal_1858, signal_1253}), .c ({DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_139 ( .a ({signal_2733, signal_2731}), .b ({signal_1859, signal_1254}), .c ({DataOut_s1[21], DataOut_s0[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_140 ( .a ({signal_2737, signal_2735}), .b ({signal_1860, signal_1255}), .c ({DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_141 ( .a ({signal_2741, signal_2739}), .b ({signal_1867, signal_1262}), .c ({DataOut_s1[1], DataOut_s0[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_142 ( .a ({signal_2745, signal_2743}), .b ({signal_1877, signal_1272}), .c ({DataOut_s1[19], DataOut_s0[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_143 ( .a ({signal_2749, signal_2747}), .b ({signal_1878, signal_1273}), .c ({DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_144 ( .a ({signal_2753, signal_2751}), .b ({signal_1879, signal_1274}), .c ({DataOut_s1[17], DataOut_s0[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_145 ( .a ({signal_2757, signal_2755}), .b ({signal_1880, signal_1275}), .c ({DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_146 ( .a ({signal_2761, signal_2759}), .b ({signal_1893, signal_1288}), .c ({DataOut_s1[15], DataOut_s0[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_147 ( .a ({signal_2765, signal_2763}), .b ({signal_1894, signal_1289}), .c ({DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_148 ( .a ({signal_2769, signal_2767}), .b ({signal_1895, signal_1290}), .c ({DataOut_s1[13], DataOut_s0[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_149 ( .a ({signal_2773, signal_2771}), .b ({signal_1896, signal_1291}), .c ({DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_150 ( .a ({signal_2777, signal_2775}), .b ({signal_1905, signal_1300}), .c ({DataOut_s1[11], DataOut_s0[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_151 ( .a ({signal_2781, signal_2779}), .b ({signal_1906, signal_1301}), .c ({DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_152 ( .a ({signal_2785, signal_2783}), .b ({signal_1868, signal_1263}), .c ({DataOut_s1[0], DataOut_s0[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_217 ( .a ({signal_2789, signal_2787}), .b ({signal_1907, signal_1302}), .c ({signal_1981, signal_1238}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_218 ( .a ({signal_1908, signal_1303}), .b ({signal_2793, signal_2791}), .c ({signal_2306, signal_1239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_219 ( .a ({signal_2797, signal_2795}), .b ({signal_1869, signal_1264}), .c ({signal_2042, signal_1240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_220 ( .a ({signal_2801, signal_2799}), .b ({signal_1870, signal_1265}), .c ({signal_2043, signal_1241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_221 ( .a ({signal_2805, signal_2803}), .b ({signal_1853, signal_1248}), .c ({signal_2044, signal_1184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_222 ( .a ({signal_2809, signal_2807}), .b ({signal_1854, signal_1249}), .c ({signal_2045, signal_1185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_223 ( .a ({signal_2813, signal_2811}), .b ({signal_1855, signal_1250}), .c ({signal_2046, signal_1186}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_224 ( .a ({signal_1856, signal_1251}), .b ({signal_2817, signal_2815}), .c ({signal_2362, signal_1187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_225 ( .a ({signal_2821, signal_2819}), .b ({signal_1871, signal_1266}), .c ({signal_2047, signal_1242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_226 ( .a ({signal_2825, signal_2823}), .b ({signal_1881, signal_1276}), .c ({signal_2048, signal_1188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_227 ( .a ({signal_2829, signal_2827}), .b ({signal_1882, signal_1277}), .c ({signal_2049, signal_1189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_228 ( .a ({signal_2833, signal_2831}), .b ({signal_1883, signal_1278}), .c ({signal_2050, signal_1190}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_229 ( .a ({signal_1884, signal_1279}), .b ({signal_2837, signal_2835}), .c ({signal_2363, signal_1191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_230 ( .a ({signal_2841, signal_2839}), .b ({signal_1909, signal_1304}), .c ({signal_2051, signal_1192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_231 ( .a ({signal_2845, signal_2843}), .b ({signal_1910, signal_1305}), .c ({signal_2052, signal_1193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_232 ( .a ({signal_2849, signal_2847}), .b ({signal_1911, signal_1306}), .c ({signal_2053, signal_1194}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_233 ( .a ({signal_1912, signal_1307}), .b ({signal_2853, signal_2851}), .c ({signal_2364, signal_1195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_234 ( .a ({signal_2857, signal_2855}), .b ({signal_1889, signal_1284}), .c ({signal_2054, signal_1196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_235 ( .a ({signal_2861, signal_2859}), .b ({signal_1890, signal_1285}), .c ({signal_2055, signal_1197}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_236 ( .a ({signal_1872, signal_1267}), .b ({signal_2865, signal_2863}), .c ({signal_2365, signal_1243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_237 ( .a ({signal_2869, signal_2867}), .b ({signal_1891, signal_1286}), .c ({signal_2056, signal_1198}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_238 ( .a ({signal_1892, signal_1287}), .b ({signal_2873, signal_2871}), .c ({signal_2389, signal_1199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_239 ( .a ({signal_2877, signal_2875}), .b ({signal_1873, signal_1268}), .c ({signal_2057, signal_1200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_240 ( .a ({signal_2881, signal_2879}), .b ({signal_1874, signal_1269}), .c ({signal_2058, signal_1201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_241 ( .a ({signal_2885, signal_2883}), .b ({signal_1875, signal_1270}), .c ({signal_2059, signal_1202}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_242 ( .a ({signal_1876, signal_1271}), .b ({signal_2889, signal_2887}), .c ({signal_2307, signal_1203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_243 ( .a ({signal_2893, signal_2891}), .b ({signal_1861, signal_1256}), .c ({signal_2060, signal_1204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_244 ( .a ({signal_2897, signal_2895}), .b ({signal_1862, signal_1257}), .c ({signal_2061, signal_1205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_245 ( .a ({signal_2901, signal_2899}), .b ({signal_1863, signal_1258}), .c ({signal_2062, signal_1206}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_246 ( .a ({signal_1864, signal_1259}), .b ({signal_2905, signal_2903}), .c ({signal_2366, signal_1207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_247 ( .a ({signal_2909, signal_2907}), .b ({signal_1865, signal_1260}), .c ({signal_1982, signal_1244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_248 ( .a ({signal_2913, signal_2911}), .b ({signal_1897, signal_1292}), .c ({signal_2063, signal_1208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_249 ( .a ({signal_2917, signal_2915}), .b ({signal_1898, signal_1293}), .c ({signal_2064, signal_1209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_250 ( .a ({signal_2921, signal_2919}), .b ({signal_1899, signal_1294}), .c ({signal_2065, signal_1210}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_251 ( .a ({signal_1900, signal_1295}), .b ({signal_2925, signal_2923}), .c ({signal_2308, signal_1211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_252 ( .a ({signal_2929, signal_2927}), .b ({signal_1901, signal_1296}), .c ({signal_2066, signal_1212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_253 ( .a ({signal_2933, signal_2931}), .b ({signal_1902, signal_1297}), .c ({signal_2067, signal_1213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_254 ( .a ({signal_2937, signal_2935}), .b ({signal_1903, signal_1298}), .c ({signal_2068, signal_1214}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_255 ( .a ({signal_1904, signal_1299}), .b ({signal_2941, signal_2939}), .c ({signal_2367, signal_1215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_256 ( .a ({signal_2945, signal_2943}), .b ({signal_1913, signal_1308}), .c ({signal_2069, signal_1216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_257 ( .a ({signal_2949, signal_2947}), .b ({signal_1914, signal_1309}), .c ({signal_2070, signal_1217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_258 ( .a ({signal_2953, signal_2951}), .b ({signal_1866, signal_1261}), .c ({signal_1983, signal_1245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_259 ( .a ({signal_2957, signal_2955}), .b ({signal_1915, signal_1310}), .c ({signal_2071, signal_1218}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_260 ( .a ({signal_1916, signal_1311}), .b ({signal_2961, signal_2959}), .c ({signal_2377, signal_1219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_261 ( .a ({signal_2965, signal_2963}), .b ({signal_1885, signal_1280}), .c ({signal_2072, signal_1220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_262 ( .a ({signal_2969, signal_2967}), .b ({signal_1886, signal_1281}), .c ({signal_1984, signal_1221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_263 ( .a ({signal_2973, signal_2971}), .b ({signal_1887, signal_1282}), .c ({signal_2073, signal_1222}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_264 ( .a ({signal_1888, signal_1283}), .b ({signal_2977, signal_2975}), .c ({signal_2368, signal_1223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_265 ( .a ({signal_2981, signal_2979}), .b ({signal_1857, signal_1252}), .c ({signal_2074, signal_1224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_266 ( .a ({signal_2985, signal_2983}), .b ({signal_1858, signal_1253}), .c ({signal_2075, signal_1225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_267 ( .a ({signal_2989, signal_2987}), .b ({signal_1859, signal_1254}), .c ({signal_2076, signal_1226}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_268 ( .a ({signal_1860, signal_1255}), .b ({signal_2993, signal_2991}), .c ({signal_2309, signal_1227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_269 ( .a ({signal_2997, signal_2995}), .b ({signal_1867, signal_1262}), .c ({signal_1985, signal_1246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_270 ( .a ({signal_3001, signal_2999}), .b ({signal_1877, signal_1272}), .c ({signal_2077, signal_1228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_271 ( .a ({signal_3005, signal_3003}), .b ({signal_1878, signal_1273}), .c ({signal_2078, signal_1229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_272 ( .a ({signal_3009, signal_3007}), .b ({signal_1879, signal_1274}), .c ({signal_2079, signal_1230}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_273 ( .a ({signal_1880, signal_1275}), .b ({signal_3013, signal_3011}), .c ({signal_2369, signal_1231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_274 ( .a ({signal_3017, signal_3015}), .b ({signal_1893, signal_1288}), .c ({signal_1986, signal_1232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_275 ( .a ({signal_3021, signal_3019}), .b ({signal_1894, signal_1289}), .c ({signal_1987, signal_1233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_276 ( .a ({signal_3025, signal_3023}), .b ({signal_1895, signal_1290}), .c ({signal_1988, signal_1234}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_277 ( .a ({signal_1896, signal_1291}), .b ({signal_3029, signal_3027}), .c ({signal_2370, signal_1235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_278 ( .a ({signal_3033, signal_3031}), .b ({signal_1905, signal_1300}), .c ({signal_1989, signal_1236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_279 ( .a ({signal_3037, signal_3035}), .b ({signal_1906, signal_1301}), .c ({signal_1990, signal_1237}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_280 ( .a ({signal_1868, signal_1263}), .b ({signal_3041, signal_3039}), .c ({signal_2371, signal_1247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_281 ( .a ({signal_2789, signal_2787}), .b ({signal_2200, signal_1110}), .c ({signal_2206, signal_1046}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_282 ( .a ({signal_2406, signal_1111}), .b ({signal_2793, signal_2791}), .c ({signal_2410, signal_1047}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_284 ( .a ({signal_2797, signal_2795}), .b ({signal_2149, signal_1064}), .c ({signal_2158, signal_1048}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_285 ( .a ({signal_2801, signal_2799}), .b ({signal_2150, signal_1065}), .c ({signal_2159, signal_1049}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_286 ( .a ({signal_2805, signal_2803}), .b ({signal_2171, signal_1056}), .c ({signal_2207, signal_992}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_287 ( .a ({signal_2809, signal_2807}), .b ({signal_2172, signal_1057}), .c ({signal_2208, signal_993}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_288 ( .a ({signal_2813, signal_2811}), .b ({signal_2173, signal_1058}), .c ({signal_2209, signal_994}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_289 ( .a ({signal_2429, signal_1059}), .b ({signal_2817, signal_2815}), .c ({signal_2441, signal_995}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_291 ( .a ({signal_2821, signal_2819}), .b ({signal_2151, signal_1066}), .c ({signal_2160, signal_1050}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_292 ( .a ({signal_2825, signal_2823}), .b ({signal_2174, signal_1096}), .c ({signal_2210, signal_996}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_293 ( .a ({signal_2829, signal_2827}), .b ({signal_2175, signal_1097}), .c ({signal_2211, signal_997}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_294 ( .a ({signal_2833, signal_2831}), .b ({signal_2164, signal_1098}), .c ({signal_2212, signal_998}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_295 ( .a ({signal_2428, signal_1099}), .b ({signal_2837, signal_2835}), .c ({signal_2442, signal_999}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_297 ( .a ({signal_2841, signal_2839}), .b ({signal_2165, signal_1076}), .c ({signal_2213, signal_1000}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_298 ( .a ({signal_2845, signal_2843}), .b ({signal_2166, signal_1077}), .c ({signal_2214, signal_1001}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_299 ( .a ({signal_2849, signal_2847}), .b ({signal_2167, signal_1078}), .c ({signal_2215, signal_1002}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_300 ( .a ({signal_2421, signal_1079}), .b ({signal_2853, signal_2851}), .c ({signal_2425, signal_1003}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_302 ( .a ({signal_2857, signal_2855}), .b ({signal_2168, signal_1116}), .c ({signal_2216, signal_1004}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_303 ( .a ({signal_2861, signal_2859}), .b ({signal_2169, signal_1117}), .c ({signal_2217, signal_1005}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_304 ( .a ({signal_2407, signal_1067}), .b ({signal_2865, signal_2863}), .c ({signal_2411, signal_1051}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_306 ( .a ({signal_2869, signal_2867}), .b ({signal_2170, signal_1118}), .c ({signal_2218, signal_1006}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_307 ( .a ({signal_2398, signal_1119}), .b ({signal_2873, signal_2871}), .c ({signal_2412, signal_1007}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_309 ( .a ({signal_2877, signal_2875}), .b ({signal_2183, signal_1112}), .c ({signal_2219, signal_1008}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_310 ( .a ({signal_2881, signal_2879}), .b ({signal_2184, signal_1113}), .c ({signal_2220, signal_1009}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_311 ( .a ({signal_2885, signal_2883}), .b ({signal_2185, signal_1114}), .c ({signal_2221, signal_1010}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_312 ( .a ({signal_2401, signal_1115}), .b ({signal_2889, signal_2887}), .c ({signal_2413, signal_1011}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_314 ( .a ({signal_2893, signal_2891}), .b ({signal_2186, signal_1072}), .c ({signal_2222, signal_1012}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_315 ( .a ({signal_2897, signal_2895}), .b ({signal_2187, signal_1073}), .c ({signal_2223, signal_1013}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_316 ( .a ({signal_2901, signal_2899}), .b ({signal_2176, signal_1074}), .c ({signal_2224, signal_1014}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_317 ( .a ({signal_2399, signal_1075}), .b ({signal_2905, signal_2903}), .c ({signal_2414, signal_1015}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_319 ( .a ({signal_2909, signal_2907}), .b ({signal_2152, signal_1088}), .c ({signal_2161, signal_1052}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_320 ( .a ({signal_2913, signal_2911}), .b ({signal_2177, signal_1100}), .c ({signal_2225, signal_1016}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_321 ( .a ({signal_2917, signal_2915}), .b ({signal_2178, signal_1101}), .c ({signal_2226, signal_1017}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_322 ( .a ({signal_2921, signal_2919}), .b ({signal_2179, signal_1102}), .c ({signal_2227, signal_1018}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_323 ( .a ({signal_2400, signal_1103}), .b ({signal_2925, signal_2923}), .c ({signal_2415, signal_1019}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_325 ( .a ({signal_2929, signal_2927}), .b ({signal_2180, signal_1060}), .c ({signal_2228, signal_1020}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_326 ( .a ({signal_2933, signal_2931}), .b ({signal_2181, signal_1061}), .c ({signal_2229, signal_1021}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_327 ( .a ({signal_2937, signal_2935}), .b ({signal_2182, signal_1062}), .c ({signal_2230, signal_1022}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_328 ( .a ({signal_2402, signal_1063}), .b ({signal_2941, signal_2939}), .c ({signal_2416, signal_1023}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_330 ( .a ({signal_2945, signal_2943}), .b ({signal_2195, signal_1092}), .c ({signal_2231, signal_1024}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_331 ( .a ({signal_2949, signal_2947}), .b ({signal_2196, signal_1093}), .c ({signal_2232, signal_1025}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_332 ( .a ({signal_2953, signal_2951}), .b ({signal_2153, signal_1089}), .c ({signal_2162, signal_1053}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_333 ( .a ({signal_2957, signal_2955}), .b ({signal_2197, signal_1094}), .c ({signal_2233, signal_1026}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_334 ( .a ({signal_2404, signal_1095}), .b ({signal_2961, signal_2959}), .c ({signal_2417, signal_1027}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_336 ( .a ({signal_2965, signal_2963}), .b ({signal_2198, signal_1068}), .c ({signal_2234, signal_1028}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_337 ( .a ({signal_2969, signal_2967}), .b ({signal_2199, signal_1069}), .c ({signal_2235, signal_1029}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_338 ( .a ({signal_2973, signal_2971}), .b ({signal_2188, signal_1070}), .c ({signal_2236, signal_1030}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_339 ( .a ({signal_2403, signal_1071}), .b ({signal_2977, signal_2975}), .c ({signal_2418, signal_1031}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_341 ( .a ({signal_2981, signal_2979}), .b ({signal_2189, signal_1104}), .c ({signal_2237, signal_1032}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_342 ( .a ({signal_2985, signal_2983}), .b ({signal_2190, signal_1105}), .c ({signal_2238, signal_1033}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_343 ( .a ({signal_2989, signal_2987}), .b ({signal_2191, signal_1106}), .c ({signal_2239, signal_1034}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_344 ( .a ({signal_2423, signal_1107}), .b ({signal_2993, signal_2991}), .c ({signal_2426, signal_1035}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_346 ( .a ({signal_2997, signal_2995}), .b ({signal_2154, signal_1090}), .c ({signal_2163, signal_1054}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_347 ( .a ({signal_3001, signal_2999}), .b ({signal_2192, signal_1080}), .c ({signal_2240, signal_1036}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_348 ( .a ({signal_3005, signal_3003}), .b ({signal_2193, signal_1081}), .c ({signal_2241, signal_1037}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_349 ( .a ({signal_3009, signal_3007}), .b ({signal_2194, signal_1082}), .c ({signal_2242, signal_1038}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_350 ( .a ({signal_2424, signal_1083}), .b ({signal_3013, signal_3011}), .c ({signal_2427, signal_1039}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_352 ( .a ({signal_3017, signal_3015}), .b ({signal_2201, signal_1084}), .c ({signal_2243, signal_1040}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_353 ( .a ({signal_3021, signal_3019}), .b ({signal_2202, signal_1085}), .c ({signal_2244, signal_1041}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_354 ( .a ({signal_3025, signal_3023}), .b ({signal_2203, signal_1086}), .c ({signal_2245, signal_1042}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_355 ( .a ({signal_2408, signal_1087}), .b ({signal_3029, signal_3027}), .c ({signal_2419, signal_1043}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_357 ( .a ({signal_3033, signal_3031}), .b ({signal_2204, signal_1108}), .c ({signal_2246, signal_1044}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_358 ( .a ({signal_3037, signal_3035}), .b ({signal_2205, signal_1109}), .c ({signal_2247, signal_1045}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_359 ( .a ({signal_2409, signal_1091}), .b ({signal_3041, signal_3039}), .c ({signal_2420, signal_1055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_535 ( .s (signal_3043), .b ({signal_2430, signal_1439}), .a ({signal_3047, signal_3045}), .c ({signal_2443, signal_460}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_538 ( .s (signal_3043), .b ({signal_2248, signal_1438}), .a ({signal_3051, signal_3049}), .c ({signal_2258, signal_462}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_541 ( .s (signal_3043), .b ({signal_2249, signal_1437}), .a ({signal_3055, signal_3053}), .c ({signal_2259, signal_464}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_544 ( .s (signal_3043), .b ({signal_2250, signal_1436}), .a ({signal_3059, signal_3057}), .c ({signal_2260, signal_466}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_547 ( .s (signal_3043), .b ({signal_2431, signal_1435}), .a ({signal_3063, signal_3061}), .c ({signal_2444, signal_468}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_550 ( .s (signal_3043), .b ({signal_2251, signal_1434}), .a ({signal_3067, signal_3065}), .c ({signal_2261, signal_470}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_553 ( .s (signal_3043), .b ({signal_2252, signal_1433}), .a ({signal_3071, signal_3069}), .c ({signal_2262, signal_472}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_556 ( .s (signal_3043), .b ({signal_2253, signal_1432}), .a ({signal_3075, signal_3073}), .c ({signal_2263, signal_474}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_559 ( .s (signal_3043), .b ({signal_2432, signal_1431}), .a ({signal_3079, signal_3077}), .c ({signal_2445, signal_476}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_562 ( .s (signal_3043), .b ({signal_2264, signal_1430}), .a ({signal_3083, signal_3081}), .c ({signal_2320, signal_478}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_565 ( .s (signal_3043), .b ({signal_2265, signal_1429}), .a ({signal_3087, signal_3085}), .c ({signal_2321, signal_480}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_568 ( .s (signal_3043), .b ({signal_2266, signal_1428}), .a ({signal_3091, signal_3089}), .c ({signal_2322, signal_482}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_571 ( .s (signal_3043), .b ({signal_2433, signal_1427}), .a ({signal_3095, signal_3093}), .c ({signal_2446, signal_484}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_574 ( .s (signal_3043), .b ({signal_2267, signal_1426}), .a ({signal_3099, signal_3097}), .c ({signal_2323, signal_486}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_577 ( .s (signal_3043), .b ({signal_2268, signal_1425}), .a ({signal_3103, signal_3101}), .c ({signal_2324, signal_488}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_580 ( .s (signal_3043), .b ({signal_2269, signal_1424}), .a ({signal_3107, signal_3105}), .c ({signal_2325, signal_490}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_583 ( .s (signal_3043), .b ({signal_2454, signal_1423}), .a ({signal_3111, signal_3109}), .c ({signal_2457, signal_492}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_586 ( .s (signal_3043), .b ({signal_2270, signal_1422}), .a ({signal_3115, signal_3113}), .c ({signal_2326, signal_494}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_589 ( .s (signal_3043), .b ({signal_2271, signal_1421}), .a ({signal_3119, signal_3117}), .c ({signal_2327, signal_496}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_592 ( .s (signal_3043), .b ({signal_2272, signal_1420}), .a ({signal_3123, signal_3121}), .c ({signal_2328, signal_498}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_595 ( .s (signal_3043), .b ({signal_2455, signal_1419}), .a ({signal_3127, signal_3125}), .c ({signal_2458, signal_500}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_598 ( .s (signal_3043), .b ({signal_2273, signal_1418}), .a ({signal_3131, signal_3129}), .c ({signal_2329, signal_502}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_601 ( .s (signal_3043), .b ({signal_2274, signal_1417}), .a ({signal_3135, signal_3133}), .c ({signal_2330, signal_504}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_604 ( .s (signal_3043), .b ({signal_2275, signal_1416}), .a ({signal_3139, signal_3137}), .c ({signal_2331, signal_506}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_607 ( .s (signal_3043), .b ({signal_2434, signal_1415}), .a ({signal_3143, signal_3141}), .c ({signal_2447, signal_508}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_610 ( .s (signal_3043), .b ({signal_2276, signal_1414}), .a ({signal_3147, signal_3145}), .c ({signal_2332, signal_510}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_613 ( .s (signal_3043), .b ({signal_2277, signal_1413}), .a ({signal_3151, signal_3149}), .c ({signal_2333, signal_512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_616 ( .s (signal_3043), .b ({signal_2278, signal_1412}), .a ({signal_3155, signal_3153}), .c ({signal_2334, signal_514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_619 ( .s (signal_3043), .b ({signal_2435, signal_1411}), .a ({signal_3159, signal_3157}), .c ({signal_2448, signal_516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_622 ( .s (signal_3043), .b ({signal_2279, signal_1410}), .a ({signal_3163, signal_3161}), .c ({signal_2335, signal_518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_625 ( .s (signal_3043), .b ({signal_2280, signal_1409}), .a ({signal_3167, signal_3165}), .c ({signal_2336, signal_520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_628 ( .s (signal_3043), .b ({signal_2281, signal_1408}), .a ({signal_3171, signal_3169}), .c ({signal_2337, signal_522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_631 ( .s (signal_3043), .b ({signal_2436, signal_1407}), .a ({signal_3175, signal_3173}), .c ({signal_2449, signal_524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_634 ( .s (signal_3043), .b ({signal_2282, signal_1406}), .a ({signal_3179, signal_3177}), .c ({signal_2338, signal_526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_637 ( .s (signal_3043), .b ({signal_2283, signal_1405}), .a ({signal_3183, signal_3181}), .c ({signal_2339, signal_528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_640 ( .s (signal_3043), .b ({signal_2284, signal_1404}), .a ({signal_3187, signal_3185}), .c ({signal_2340, signal_530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_643 ( .s (signal_3043), .b ({signal_2437, signal_1403}), .a ({signal_3191, signal_3189}), .c ({signal_2450, signal_532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_646 ( .s (signal_3043), .b ({signal_2285, signal_1402}), .a ({signal_3195, signal_3193}), .c ({signal_2341, signal_534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_649 ( .s (signal_3043), .b ({signal_2286, signal_1401}), .a ({signal_3199, signal_3197}), .c ({signal_2342, signal_536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_652 ( .s (signal_3043), .b ({signal_2287, signal_1400}), .a ({signal_3203, signal_3201}), .c ({signal_2343, signal_538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_655 ( .s (signal_3043), .b ({signal_2438, signal_1399}), .a ({signal_3207, signal_3205}), .c ({signal_2451, signal_540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_658 ( .s (signal_3043), .b ({signal_2288, signal_1398}), .a ({signal_3211, signal_3209}), .c ({signal_2344, signal_542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_661 ( .s (signal_3043), .b ({signal_2289, signal_1397}), .a ({signal_3215, signal_3213}), .c ({signal_2345, signal_544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_664 ( .s (signal_3043), .b ({signal_2290, signal_1396}), .a ({signal_3219, signal_3217}), .c ({signal_2346, signal_546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_667 ( .s (signal_3043), .b ({signal_2439, signal_1395}), .a ({signal_3223, signal_3221}), .c ({signal_2452, signal_548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_670 ( .s (signal_3043), .b ({signal_2291, signal_1394}), .a ({signal_3227, signal_3225}), .c ({signal_2347, signal_550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_673 ( .s (signal_3043), .b ({signal_2292, signal_1393}), .a ({signal_3231, signal_3229}), .c ({signal_2348, signal_552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_676 ( .s (signal_3043), .b ({signal_2293, signal_1392}), .a ({signal_3235, signal_3233}), .c ({signal_2349, signal_554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_679 ( .s (signal_3043), .b ({signal_2440, signal_1391}), .a ({signal_3239, signal_3237}), .c ({signal_2453, signal_556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_682 ( .s (signal_3043), .b ({signal_2294, signal_1390}), .a ({signal_3243, signal_3241}), .c ({signal_2350, signal_558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_685 ( .s (signal_3043), .b ({signal_2295, signal_1389}), .a ({signal_3247, signal_3245}), .c ({signal_2351, signal_560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_688 ( .s (signal_3043), .b ({signal_2296, signal_1388}), .a ({signal_3251, signal_3249}), .c ({signal_2352, signal_562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_691 ( .s (signal_3043), .b ({signal_2456, signal_1387}), .a ({signal_3255, signal_3253}), .c ({signal_2459, signal_564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_694 ( .s (signal_3043), .b ({signal_2297, signal_1386}), .a ({signal_3259, signal_3257}), .c ({signal_2353, signal_566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_697 ( .s (signal_3043), .b ({signal_2298, signal_1385}), .a ({signal_3263, signal_3261}), .c ({signal_2354, signal_568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_700 ( .s (signal_3043), .b ({signal_2299, signal_1384}), .a ({signal_3267, signal_3265}), .c ({signal_2355, signal_570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_703 ( .s (signal_3043), .b ({signal_2460, signal_1383}), .a ({signal_3271, signal_3269}), .c ({signal_2462, signal_572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_706 ( .s (signal_3043), .b ({signal_2300, signal_1382}), .a ({signal_3275, signal_3273}), .c ({signal_2356, signal_574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_709 ( .s (signal_3043), .b ({signal_2301, signal_1381}), .a ({signal_3279, signal_3277}), .c ({signal_2357, signal_576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_712 ( .s (signal_3043), .b ({signal_2302, signal_1380}), .a ({signal_3283, signal_3281}), .c ({signal_2358, signal_578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_715 ( .s (signal_3043), .b ({signal_2461, signal_1379}), .a ({signal_3287, signal_3285}), .c ({signal_2463, signal_580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_718 ( .s (signal_3043), .b ({signal_2303, signal_1378}), .a ({signal_3291, signal_3289}), .c ({signal_2359, signal_582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_721 ( .s (signal_3043), .b ({signal_2304, signal_1377}), .a ({signal_3295, signal_3293}), .c ({signal_2360, signal_584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_724 ( .s (signal_3043), .b ({signal_2305, signal_1376}), .a ({signal_3299, signal_3297}), .c ({signal_2361, signal_586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1031 ( .s (signal_3301), .b ({signal_1916, signal_1311}), .a ({signal_2371, signal_1247}), .c ({signal_2379, signal_1183}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1032 ( .s (signal_3301), .b ({signal_1915, signal_1310}), .a ({signal_1985, signal_1246}), .c ({signal_2080, signal_1182}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1033 ( .s (signal_3301), .b ({signal_1914, signal_1309}), .a ({signal_1983, signal_1245}), .c ({signal_2081, signal_1181}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1034 ( .s (signal_3301), .b ({signal_1913, signal_1308}), .a ({signal_1982, signal_1244}), .c ({signal_2082, signal_1180}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1035 ( .s (signal_3301), .b ({signal_1912, signal_1307}), .a ({signal_2365, signal_1243}), .c ({signal_2380, signal_1179}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1036 ( .s (signal_3301), .b ({signal_1911, signal_1306}), .a ({signal_2047, signal_1242}), .c ({signal_2090, signal_1178}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1037 ( .s (signal_3301), .b ({signal_1910, signal_1305}), .a ({signal_2043, signal_1241}), .c ({signal_2091, signal_1177}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1038 ( .s (signal_3301), .b ({signal_1909, signal_1304}), .a ({signal_2042, signal_1240}), .c ({signal_2092, signal_1176}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1039 ( .s (signal_3301), .b ({signal_1908, signal_1303}), .a ({signal_2306, signal_1239}), .c ({signal_2373, signal_1175}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1040 ( .s (signal_3301), .b ({signal_1907, signal_1302}), .a ({signal_1981, signal_1238}), .c ({signal_2083, signal_1174}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1041 ( .s (signal_3301), .b ({signal_1906, signal_1301}), .a ({signal_1990, signal_1237}), .c ({signal_2084, signal_1173}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1042 ( .s (signal_3301), .b ({signal_1905, signal_1300}), .a ({signal_1989, signal_1236}), .c ({signal_2085, signal_1172}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1043 ( .s (signal_3301), .b ({signal_1904, signal_1299}), .a ({signal_2370, signal_1235}), .c ({signal_2381, signal_1171}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1044 ( .s (signal_3301), .b ({signal_1903, signal_1298}), .a ({signal_1988, signal_1234}), .c ({signal_2086, signal_1170}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1045 ( .s (signal_3301), .b ({signal_1902, signal_1297}), .a ({signal_1987, signal_1233}), .c ({signal_2087, signal_1169}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1046 ( .s (signal_3301), .b ({signal_1901, signal_1296}), .a ({signal_1986, signal_1232}), .c ({signal_2088, signal_1168}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1047 ( .s (signal_3301), .b ({signal_1900, signal_1295}), .a ({signal_2369, signal_1231}), .c ({signal_2382, signal_1167}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1048 ( .s (signal_3301), .b ({signal_1899, signal_1294}), .a ({signal_2079, signal_1230}), .c ({signal_2093, signal_1166}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1049 ( .s (signal_3301), .b ({signal_1898, signal_1293}), .a ({signal_2078, signal_1229}), .c ({signal_2094, signal_1165}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1050 ( .s (signal_3301), .b ({signal_1897, signal_1292}), .a ({signal_2077, signal_1228}), .c ({signal_2095, signal_1164}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1051 ( .s (signal_3301), .b ({signal_1896, signal_1291}), .a ({signal_2309, signal_1227}), .c ({signal_2374, signal_1163}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1052 ( .s (signal_3301), .b ({signal_1895, signal_1290}), .a ({signal_2076, signal_1226}), .c ({signal_2096, signal_1162}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1053 ( .s (signal_3301), .b ({signal_1894, signal_1289}), .a ({signal_2075, signal_1225}), .c ({signal_2097, signal_1161}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1054 ( .s (signal_3301), .b ({signal_1893, signal_1288}), .a ({signal_2074, signal_1224}), .c ({signal_2098, signal_1160}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1055 ( .s (signal_3301), .b ({signal_1892, signal_1287}), .a ({signal_2368, signal_1223}), .c ({signal_2383, signal_1159}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1056 ( .s (signal_3301), .b ({signal_1891, signal_1286}), .a ({signal_2073, signal_1222}), .c ({signal_2099, signal_1158}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1057 ( .s (signal_3301), .b ({signal_1890, signal_1285}), .a ({signal_1984, signal_1221}), .c ({signal_2089, signal_1157}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1058 ( .s (signal_3301), .b ({signal_1889, signal_1284}), .a ({signal_2072, signal_1220}), .c ({signal_2100, signal_1156}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1059 ( .s (signal_3301), .b ({signal_1888, signal_1283}), .a ({signal_2377, signal_1219}), .c ({signal_2390, signal_1155}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1060 ( .s (signal_3301), .b ({signal_1887, signal_1282}), .a ({signal_2071, signal_1218}), .c ({signal_2101, signal_1154}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1061 ( .s (signal_3301), .b ({signal_1886, signal_1281}), .a ({signal_2070, signal_1217}), .c ({signal_2102, signal_1153}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1062 ( .s (signal_3301), .b ({signal_1885, signal_1280}), .a ({signal_2069, signal_1216}), .c ({signal_2103, signal_1152}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1063 ( .s (signal_3301), .b ({signal_1884, signal_1279}), .a ({signal_2367, signal_1215}), .c ({signal_2384, signal_1151}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1064 ( .s (signal_3301), .b ({signal_1883, signal_1278}), .a ({signal_2068, signal_1214}), .c ({signal_2104, signal_1150}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1065 ( .s (signal_3301), .b ({signal_1882, signal_1277}), .a ({signal_2067, signal_1213}), .c ({signal_2105, signal_1149}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1066 ( .s (signal_3301), .b ({signal_1881, signal_1276}), .a ({signal_2066, signal_1212}), .c ({signal_2106, signal_1148}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1067 ( .s (signal_3301), .b ({signal_1880, signal_1275}), .a ({signal_2308, signal_1211}), .c ({signal_2375, signal_1147}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1068 ( .s (signal_3301), .b ({signal_1879, signal_1274}), .a ({signal_2065, signal_1210}), .c ({signal_2107, signal_1146}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1069 ( .s (signal_3301), .b ({signal_1878, signal_1273}), .a ({signal_2064, signal_1209}), .c ({signal_2108, signal_1145}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1070 ( .s (signal_3301), .b ({signal_1877, signal_1272}), .a ({signal_2063, signal_1208}), .c ({signal_2109, signal_1144}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1071 ( .s (signal_3301), .b ({signal_1876, signal_1271}), .a ({signal_2366, signal_1207}), .c ({signal_2385, signal_1143}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1072 ( .s (signal_3301), .b ({signal_1875, signal_1270}), .a ({signal_2062, signal_1206}), .c ({signal_2110, signal_1142}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1073 ( .s (signal_3301), .b ({signal_1874, signal_1269}), .a ({signal_2061, signal_1205}), .c ({signal_2111, signal_1141}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1074 ( .s (signal_3301), .b ({signal_1873, signal_1268}), .a ({signal_2060, signal_1204}), .c ({signal_2112, signal_1140}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1075 ( .s (signal_3301), .b ({signal_1872, signal_1267}), .a ({signal_2307, signal_1203}), .c ({signal_2376, signal_1139}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1076 ( .s (signal_3301), .b ({signal_1871, signal_1266}), .a ({signal_2059, signal_1202}), .c ({signal_2113, signal_1138}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1077 ( .s (signal_3301), .b ({signal_1870, signal_1265}), .a ({signal_2058, signal_1201}), .c ({signal_2114, signal_1137}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1078 ( .s (signal_3301), .b ({signal_1869, signal_1264}), .a ({signal_2057, signal_1200}), .c ({signal_2115, signal_1136}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1079 ( .s (signal_3301), .b ({signal_1868, signal_1263}), .a ({signal_2389, signal_1199}), .c ({signal_2397, signal_1135}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1080 ( .s (signal_3301), .b ({signal_1867, signal_1262}), .a ({signal_2056, signal_1198}), .c ({signal_2116, signal_1134}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1081 ( .s (signal_3301), .b ({signal_1866, signal_1261}), .a ({signal_2055, signal_1197}), .c ({signal_2117, signal_1133}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1082 ( .s (signal_3301), .b ({signal_1865, signal_1260}), .a ({signal_2054, signal_1196}), .c ({signal_2118, signal_1132}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1083 ( .s (signal_3301), .b ({signal_1864, signal_1259}), .a ({signal_2364, signal_1195}), .c ({signal_2386, signal_1131}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1084 ( .s (signal_3301), .b ({signal_1863, signal_1258}), .a ({signal_2053, signal_1194}), .c ({signal_2119, signal_1130}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1085 ( .s (signal_3301), .b ({signal_1862, signal_1257}), .a ({signal_2052, signal_1193}), .c ({signal_2120, signal_1129}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1086 ( .s (signal_3301), .b ({signal_1861, signal_1256}), .a ({signal_2051, signal_1192}), .c ({signal_2121, signal_1128}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1087 ( .s (signal_3301), .b ({signal_1860, signal_1255}), .a ({signal_2363, signal_1191}), .c ({signal_2387, signal_1127}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1088 ( .s (signal_3301), .b ({signal_1859, signal_1254}), .a ({signal_2050, signal_1190}), .c ({signal_2122, signal_1126}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1089 ( .s (signal_3301), .b ({signal_1858, signal_1253}), .a ({signal_2049, signal_1189}), .c ({signal_2123, signal_1125}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1090 ( .s (signal_3301), .b ({signal_1857, signal_1252}), .a ({signal_2048, signal_1188}), .c ({signal_2124, signal_1124}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1091 ( .s (signal_3301), .b ({signal_1856, signal_1251}), .a ({signal_2362, signal_1187}), .c ({signal_2388, signal_1123}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1092 ( .s (signal_3301), .b ({signal_1855, signal_1250}), .a ({signal_2046, signal_1186}), .c ({signal_2125, signal_1122}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1093 ( .s (signal_3301), .b ({signal_1854, signal_1249}), .a ({signal_2045, signal_1185}), .c ({signal_2126, signal_1121}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1094 ( .s (signal_3301), .b ({signal_1853, signal_1248}), .a ({signal_2044, signal_1184}), .c ({signal_2127, signal_1120}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1095 ( .a ({signal_2125, signal_1122}), .b ({signal_2134, signal_828}), .c ({signal_2164, signal_1098}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1096 ( .a ({signal_2388, signal_1123}), .b ({signal_2422, signal_829}), .c ({signal_2428, signal_1099}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1097 ( .a ({signal_2118, signal_1132}), .b ({signal_2131, signal_830}), .c ({signal_2165, signal_1076}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1098 ( .a ({signal_2117, signal_1133}), .b ({signal_2132, signal_831}), .c ({signal_2166, signal_1077}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1099 ( .a ({signal_2116, signal_1134}), .b ({signal_2133, signal_832}), .c ({signal_2167, signal_1078}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1100 ( .a ({signal_2397, signal_1135}), .b ({signal_2391, signal_833}), .c ({signal_2421, signal_1079}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1101 ( .a ({signal_2121, signal_1128}), .b ({signal_2131, signal_830}), .c ({signal_2168, signal_1116}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1102 ( .a ({signal_2127, signal_1120}), .b ({signal_2124, signal_1124}), .c ({signal_2131, signal_830}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1103 ( .a ({signal_2120, signal_1129}), .b ({signal_2132, signal_831}), .c ({signal_2169, signal_1117}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1104 ( .a ({signal_2126, signal_1121}), .b ({signal_2123, signal_1125}), .c ({signal_2132, signal_831}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1105 ( .a ({signal_2119, signal_1130}), .b ({signal_2133, signal_832}), .c ({signal_2170, signal_1118}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1106 ( .a ({signal_2122, signal_1126}), .b ({signal_2125, signal_1122}), .c ({signal_2133, signal_832}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1107 ( .a ({signal_2124, signal_1124}), .b ({signal_2135, signal_834}), .c ({signal_2171, signal_1056}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1108 ( .a ({signal_2123, signal_1125}), .b ({signal_2136, signal_835}), .c ({signal_2172, signal_1057}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1109 ( .a ({signal_2122, signal_1126}), .b ({signal_2134, signal_828}), .c ({signal_2173, signal_1058}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1110 ( .a ({signal_2116, signal_1134}), .b ({signal_2119, signal_1130}), .c ({signal_2134, signal_828}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1111 ( .a ({signal_2387, signal_1127}), .b ({signal_2422, signal_829}), .c ({signal_2429, signal_1059}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1112 ( .a ({signal_2386, signal_1131}), .b ({signal_2397, signal_1135}), .c ({signal_2422, signal_829}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1113 ( .a ({signal_2127, signal_1120}), .b ({signal_2135, signal_834}), .c ({signal_2174, signal_1096}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1114 ( .a ({signal_2118, signal_1132}), .b ({signal_2121, signal_1128}), .c ({signal_2135, signal_834}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1115 ( .a ({signal_2126, signal_1121}), .b ({signal_2136, signal_835}), .c ({signal_2175, signal_1097}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1116 ( .a ({signal_2117, signal_1133}), .b ({signal_2120, signal_1129}), .c ({signal_2136, signal_835}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1117 ( .a ({signal_2386, signal_1131}), .b ({signal_2391, signal_833}), .c ({signal_2398, signal_1119}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1118 ( .a ({signal_2388, signal_1123}), .b ({signal_2387, signal_1127}), .c ({signal_2391, signal_833}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1119 ( .a ({signal_2113, signal_1138}), .b ({signal_2140, signal_836}), .c ({signal_2176, signal_1074}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1120 ( .a ({signal_2376, signal_1139}), .b ({signal_2392, signal_837}), .c ({signal_2399, signal_1075}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1121 ( .a ({signal_2106, signal_1148}), .b ({signal_2137, signal_838}), .c ({signal_2177, signal_1100}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1122 ( .a ({signal_2105, signal_1149}), .b ({signal_2138, signal_839}), .c ({signal_2178, signal_1101}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1123 ( .a ({signal_2104, signal_1150}), .b ({signal_2139, signal_840}), .c ({signal_2179, signal_1102}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1124 ( .a ({signal_2384, signal_1151}), .b ({signal_2393, signal_841}), .c ({signal_2400, signal_1103}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1125 ( .a ({signal_2109, signal_1144}), .b ({signal_2137, signal_838}), .c ({signal_2180, signal_1060}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1126 ( .a ({signal_2115, signal_1136}), .b ({signal_2112, signal_1140}), .c ({signal_2137, signal_838}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1127 ( .a ({signal_2108, signal_1145}), .b ({signal_2138, signal_839}), .c ({signal_2181, signal_1061}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1128 ( .a ({signal_2114, signal_1137}), .b ({signal_2111, signal_1141}), .c ({signal_2138, signal_839}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1129 ( .a ({signal_2107, signal_1146}), .b ({signal_2139, signal_840}), .c ({signal_2182, signal_1062}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1130 ( .a ({signal_2110, signal_1142}), .b ({signal_2113, signal_1138}), .c ({signal_2139, signal_840}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1131 ( .a ({signal_2112, signal_1140}), .b ({signal_2141, signal_842}), .c ({signal_2183, signal_1112}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1132 ( .a ({signal_2111, signal_1141}), .b ({signal_2142, signal_843}), .c ({signal_2184, signal_1113}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1133 ( .a ({signal_2110, signal_1142}), .b ({signal_2140, signal_836}), .c ({signal_2185, signal_1114}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1134 ( .a ({signal_2104, signal_1150}), .b ({signal_2107, signal_1146}), .c ({signal_2140, signal_836}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1135 ( .a ({signal_2385, signal_1143}), .b ({signal_2392, signal_837}), .c ({signal_2401, signal_1115}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1136 ( .a ({signal_2375, signal_1147}), .b ({signal_2384, signal_1151}), .c ({signal_2392, signal_837}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1137 ( .a ({signal_2115, signal_1136}), .b ({signal_2141, signal_842}), .c ({signal_2186, signal_1072}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1138 ( .a ({signal_2106, signal_1148}), .b ({signal_2109, signal_1144}), .c ({signal_2141, signal_842}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1139 ( .a ({signal_2114, signal_1137}), .b ({signal_2142, signal_843}), .c ({signal_2187, signal_1073}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1140 ( .a ({signal_2105, signal_1149}), .b ({signal_2108, signal_1145}), .c ({signal_2142, signal_843}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1141 ( .a ({signal_2375, signal_1147}), .b ({signal_2393, signal_841}), .c ({signal_2402, signal_1063}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1142 ( .a ({signal_2376, signal_1139}), .b ({signal_2385, signal_1143}), .c ({signal_2393, signal_841}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1143 ( .a ({signal_2101, signal_1154}), .b ({signal_2146, signal_844}), .c ({signal_2188, signal_1070}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1144 ( .a ({signal_2390, signal_1155}), .b ({signal_2394, signal_845}), .c ({signal_2403, signal_1071}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1145 ( .a ({signal_2095, signal_1164}), .b ({signal_2143, signal_846}), .c ({signal_2189, signal_1104}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1146 ( .a ({signal_2094, signal_1165}), .b ({signal_2144, signal_847}), .c ({signal_2190, signal_1105}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1147 ( .a ({signal_2093, signal_1166}), .b ({signal_2145, signal_848}), .c ({signal_2191, signal_1106}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1148 ( .a ({signal_2382, signal_1167}), .b ({signal_2405, signal_849}), .c ({signal_2423, signal_1107}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1149 ( .a ({signal_2098, signal_1160}), .b ({signal_2143, signal_846}), .c ({signal_2192, signal_1080}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1150 ( .a ({signal_2103, signal_1152}), .b ({signal_2100, signal_1156}), .c ({signal_2143, signal_846}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1151 ( .a ({signal_2097, signal_1161}), .b ({signal_2144, signal_847}), .c ({signal_2193, signal_1081}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1152 ( .a ({signal_2102, signal_1153}), .b ({signal_2089, signal_1157}), .c ({signal_2144, signal_847}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1153 ( .a ({signal_2096, signal_1162}), .b ({signal_2145, signal_848}), .c ({signal_2194, signal_1082}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1154 ( .a ({signal_2099, signal_1158}), .b ({signal_2101, signal_1154}), .c ({signal_2145, signal_848}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1155 ( .a ({signal_2100, signal_1156}), .b ({signal_2147, signal_850}), .c ({signal_2195, signal_1092}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1156 ( .a ({signal_2089, signal_1157}), .b ({signal_2148, signal_851}), .c ({signal_2196, signal_1093}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1157 ( .a ({signal_2099, signal_1158}), .b ({signal_2146, signal_844}), .c ({signal_2197, signal_1094}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1158 ( .a ({signal_2093, signal_1166}), .b ({signal_2096, signal_1162}), .c ({signal_2146, signal_844}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1159 ( .a ({signal_2383, signal_1159}), .b ({signal_2394, signal_845}), .c ({signal_2404, signal_1095}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1160 ( .a ({signal_2374, signal_1163}), .b ({signal_2382, signal_1167}), .c ({signal_2394, signal_845}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1161 ( .a ({signal_2103, signal_1152}), .b ({signal_2147, signal_850}), .c ({signal_2198, signal_1068}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1162 ( .a ({signal_2095, signal_1164}), .b ({signal_2098, signal_1160}), .c ({signal_2147, signal_850}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1163 ( .a ({signal_2102, signal_1153}), .b ({signal_2148, signal_851}), .c ({signal_2199, signal_1069}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1164 ( .a ({signal_2094, signal_1165}), .b ({signal_2097, signal_1161}), .c ({signal_2148, signal_851}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1165 ( .a ({signal_2374, signal_1163}), .b ({signal_2405, signal_849}), .c ({signal_2424, signal_1083}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1166 ( .a ({signal_2390, signal_1155}), .b ({signal_2383, signal_1159}), .c ({signal_2405, signal_849}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1167 ( .a ({signal_2086, signal_1170}), .b ({signal_2155, signal_852}), .c ({signal_2200, signal_1110}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1168 ( .a ({signal_2381, signal_1171}), .b ({signal_2395, signal_853}), .c ({signal_2406, signal_1111}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1169 ( .a ({signal_2082, signal_1180}), .b ({signal_2128, signal_854}), .c ({signal_2149, signal_1064}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1170 ( .a ({signal_2081, signal_1181}), .b ({signal_2129, signal_855}), .c ({signal_2150, signal_1065}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1171 ( .a ({signal_2080, signal_1182}), .b ({signal_2130, signal_856}), .c ({signal_2151, signal_1066}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1172 ( .a ({signal_2379, signal_1183}), .b ({signal_2396, signal_857}), .c ({signal_2407, signal_1067}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1173 ( .a ({signal_2092, signal_1176}), .b ({signal_2128, signal_854}), .c ({signal_2152, signal_1088}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1174 ( .a ({signal_2088, signal_1168}), .b ({signal_2085, signal_1172}), .c ({signal_2128, signal_854}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1175 ( .a ({signal_2091, signal_1177}), .b ({signal_2129, signal_855}), .c ({signal_2153, signal_1089}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1176 ( .a ({signal_2087, signal_1169}), .b ({signal_2084, signal_1173}), .c ({signal_2129, signal_855}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1177 ( .a ({signal_2090, signal_1178}), .b ({signal_2130, signal_856}), .c ({signal_2154, signal_1090}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1178 ( .a ({signal_2083, signal_1174}), .b ({signal_2086, signal_1170}), .c ({signal_2130, signal_856}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1179 ( .a ({signal_2085, signal_1172}), .b ({signal_2156, signal_858}), .c ({signal_2201, signal_1084}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1180 ( .a ({signal_2084, signal_1173}), .b ({signal_2157, signal_859}), .c ({signal_2202, signal_1085}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1181 ( .a ({signal_2083, signal_1174}), .b ({signal_2155, signal_852}), .c ({signal_2203, signal_1086}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1182 ( .a ({signal_2080, signal_1182}), .b ({signal_2090, signal_1178}), .c ({signal_2155, signal_852}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1183 ( .a ({signal_2373, signal_1175}), .b ({signal_2395, signal_853}), .c ({signal_2408, signal_1087}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1184 ( .a ({signal_2380, signal_1179}), .b ({signal_2379, signal_1183}), .c ({signal_2395, signal_853}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1185 ( .a ({signal_2088, signal_1168}), .b ({signal_2156, signal_858}), .c ({signal_2204, signal_1108}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1186 ( .a ({signal_2082, signal_1180}), .b ({signal_2092, signal_1176}), .c ({signal_2156, signal_858}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1187 ( .a ({signal_2087, signal_1169}), .b ({signal_2157, signal_859}), .c ({signal_2205, signal_1109}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1188 ( .a ({signal_2081, signal_1181}), .b ({signal_2091, signal_1177}), .c ({signal_2157, signal_859}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1189 ( .a ({signal_2380, signal_1179}), .b ({signal_2396, signal_857}), .c ({signal_2409, signal_1091}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1190 ( .a ({signal_2381, signal_1171}), .b ({signal_2373, signal_1175}), .c ({signal_2396, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1191 ( .s (signal_3301), .b ({signal_2420, signal_1055}), .a ({signal_2398, signal_1119}), .c ({signal_2430, signal_1439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1192 ( .s (signal_3301), .b ({signal_2163, signal_1054}), .a ({signal_2170, signal_1118}), .c ({signal_2248, signal_1438}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1193 ( .s (signal_3301), .b ({signal_2162, signal_1053}), .a ({signal_2169, signal_1117}), .c ({signal_2249, signal_1437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1194 ( .s (signal_3301), .b ({signal_2161, signal_1052}), .a ({signal_2168, signal_1116}), .c ({signal_2250, signal_1436}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1195 ( .s (signal_3301), .b ({signal_2411, signal_1051}), .a ({signal_2401, signal_1115}), .c ({signal_2431, signal_1435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1196 ( .s (signal_3301), .b ({signal_2160, signal_1050}), .a ({signal_2185, signal_1114}), .c ({signal_2251, signal_1434}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1197 ( .s (signal_3301), .b ({signal_2159, signal_1049}), .a ({signal_2184, signal_1113}), .c ({signal_2252, signal_1433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1198 ( .s (signal_3301), .b ({signal_2158, signal_1048}), .a ({signal_2183, signal_1112}), .c ({signal_2253, signal_1432}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1199 ( .s (signal_3301), .b ({signal_2410, signal_1047}), .a ({signal_2406, signal_1111}), .c ({signal_2432, signal_1431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1200 ( .s (signal_3301), .b ({signal_2206, signal_1046}), .a ({signal_2200, signal_1110}), .c ({signal_2264, signal_1430}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1201 ( .s (signal_3301), .b ({signal_2247, signal_1045}), .a ({signal_2205, signal_1109}), .c ({signal_2265, signal_1429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1202 ( .s (signal_3301), .b ({signal_2246, signal_1044}), .a ({signal_2204, signal_1108}), .c ({signal_2266, signal_1428}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1203 ( .s (signal_3301), .b ({signal_2419, signal_1043}), .a ({signal_2423, signal_1107}), .c ({signal_2433, signal_1427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1204 ( .s (signal_3301), .b ({signal_2245, signal_1042}), .a ({signal_2191, signal_1106}), .c ({signal_2267, signal_1426}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1205 ( .s (signal_3301), .b ({signal_2244, signal_1041}), .a ({signal_2190, signal_1105}), .c ({signal_2268, signal_1425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1206 ( .s (signal_3301), .b ({signal_2243, signal_1040}), .a ({signal_2189, signal_1104}), .c ({signal_2269, signal_1424}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1207 ( .s (signal_3301), .b ({signal_2427, signal_1039}), .a ({signal_2400, signal_1103}), .c ({signal_2454, signal_1423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1208 ( .s (signal_3301), .b ({signal_2242, signal_1038}), .a ({signal_2179, signal_1102}), .c ({signal_2270, signal_1422}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1209 ( .s (signal_3301), .b ({signal_2241, signal_1037}), .a ({signal_2178, signal_1101}), .c ({signal_2271, signal_1421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1210 ( .s (signal_3301), .b ({signal_2240, signal_1036}), .a ({signal_2177, signal_1100}), .c ({signal_2272, signal_1420}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1211 ( .s (signal_3301), .b ({signal_2426, signal_1035}), .a ({signal_2428, signal_1099}), .c ({signal_2455, signal_1419}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1212 ( .s (signal_3301), .b ({signal_2239, signal_1034}), .a ({signal_2164, signal_1098}), .c ({signal_2273, signal_1418}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1213 ( .s (signal_3301), .b ({signal_2238, signal_1033}), .a ({signal_2175, signal_1097}), .c ({signal_2274, signal_1417}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1214 ( .s (signal_3301), .b ({signal_2237, signal_1032}), .a ({signal_2174, signal_1096}), .c ({signal_2275, signal_1416}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1215 ( .s (signal_3301), .b ({signal_2418, signal_1031}), .a ({signal_2404, signal_1095}), .c ({signal_2434, signal_1415}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1216 ( .s (signal_3301), .b ({signal_2236, signal_1030}), .a ({signal_2197, signal_1094}), .c ({signal_2276, signal_1414}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1217 ( .s (signal_3301), .b ({signal_2235, signal_1029}), .a ({signal_2196, signal_1093}), .c ({signal_2277, signal_1413}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1218 ( .s (signal_3301), .b ({signal_2234, signal_1028}), .a ({signal_2195, signal_1092}), .c ({signal_2278, signal_1412}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1219 ( .s (signal_3301), .b ({signal_2417, signal_1027}), .a ({signal_2409, signal_1091}), .c ({signal_2435, signal_1411}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1220 ( .s (signal_3301), .b ({signal_2233, signal_1026}), .a ({signal_2154, signal_1090}), .c ({signal_2279, signal_1410}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1221 ( .s (signal_3301), .b ({signal_2232, signal_1025}), .a ({signal_2153, signal_1089}), .c ({signal_2280, signal_1409}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1222 ( .s (signal_3301), .b ({signal_2231, signal_1024}), .a ({signal_2152, signal_1088}), .c ({signal_2281, signal_1408}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1223 ( .s (signal_3301), .b ({signal_2416, signal_1023}), .a ({signal_2408, signal_1087}), .c ({signal_2436, signal_1407}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1224 ( .s (signal_3301), .b ({signal_2230, signal_1022}), .a ({signal_2203, signal_1086}), .c ({signal_2282, signal_1406}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1225 ( .s (signal_3301), .b ({signal_2229, signal_1021}), .a ({signal_2202, signal_1085}), .c ({signal_2283, signal_1405}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1226 ( .s (signal_3301), .b ({signal_2228, signal_1020}), .a ({signal_2201, signal_1084}), .c ({signal_2284, signal_1404}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1227 ( .s (signal_3301), .b ({signal_2415, signal_1019}), .a ({signal_2424, signal_1083}), .c ({signal_2437, signal_1403}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1228 ( .s (signal_3301), .b ({signal_2227, signal_1018}), .a ({signal_2194, signal_1082}), .c ({signal_2285, signal_1402}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1229 ( .s (signal_3301), .b ({signal_2226, signal_1017}), .a ({signal_2193, signal_1081}), .c ({signal_2286, signal_1401}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1230 ( .s (signal_3301), .b ({signal_2225, signal_1016}), .a ({signal_2192, signal_1080}), .c ({signal_2287, signal_1400}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1231 ( .s (signal_3301), .b ({signal_2414, signal_1015}), .a ({signal_2421, signal_1079}), .c ({signal_2438, signal_1399}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1232 ( .s (signal_3301), .b ({signal_2224, signal_1014}), .a ({signal_2167, signal_1078}), .c ({signal_2288, signal_1398}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1233 ( .s (signal_3301), .b ({signal_2223, signal_1013}), .a ({signal_2166, signal_1077}), .c ({signal_2289, signal_1397}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1234 ( .s (signal_3301), .b ({signal_2222, signal_1012}), .a ({signal_2165, signal_1076}), .c ({signal_2290, signal_1396}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1235 ( .s (signal_3301), .b ({signal_2413, signal_1011}), .a ({signal_2399, signal_1075}), .c ({signal_2439, signal_1395}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1236 ( .s (signal_3301), .b ({signal_2221, signal_1010}), .a ({signal_2176, signal_1074}), .c ({signal_2291, signal_1394}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1237 ( .s (signal_3301), .b ({signal_2220, signal_1009}), .a ({signal_2187, signal_1073}), .c ({signal_2292, signal_1393}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1238 ( .s (signal_3301), .b ({signal_2219, signal_1008}), .a ({signal_2186, signal_1072}), .c ({signal_2293, signal_1392}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1239 ( .s (signal_3301), .b ({signal_2412, signal_1007}), .a ({signal_2403, signal_1071}), .c ({signal_2440, signal_1391}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1240 ( .s (signal_3301), .b ({signal_2218, signal_1006}), .a ({signal_2188, signal_1070}), .c ({signal_2294, signal_1390}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1241 ( .s (signal_3301), .b ({signal_2217, signal_1005}), .a ({signal_2199, signal_1069}), .c ({signal_2295, signal_1389}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1242 ( .s (signal_3301), .b ({signal_2216, signal_1004}), .a ({signal_2198, signal_1068}), .c ({signal_2296, signal_1388}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1243 ( .s (signal_3301), .b ({signal_2425, signal_1003}), .a ({signal_2407, signal_1067}), .c ({signal_2456, signal_1387}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1244 ( .s (signal_3301), .b ({signal_2215, signal_1002}), .a ({signal_2151, signal_1066}), .c ({signal_2297, signal_1386}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1245 ( .s (signal_3301), .b ({signal_2214, signal_1001}), .a ({signal_2150, signal_1065}), .c ({signal_2298, signal_1385}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1246 ( .s (signal_3301), .b ({signal_2213, signal_1000}), .a ({signal_2149, signal_1064}), .c ({signal_2299, signal_1384}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1247 ( .s (signal_3301), .b ({signal_2442, signal_999}), .a ({signal_2402, signal_1063}), .c ({signal_2460, signal_1383}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1248 ( .s (signal_3301), .b ({signal_2212, signal_998}), .a ({signal_2182, signal_1062}), .c ({signal_2300, signal_1382}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1249 ( .s (signal_3301), .b ({signal_2211, signal_997}), .a ({signal_2181, signal_1061}), .c ({signal_2301, signal_1381}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1250 ( .s (signal_3301), .b ({signal_2210, signal_996}), .a ({signal_2180, signal_1060}), .c ({signal_2302, signal_1380}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1251 ( .s (signal_3301), .b ({signal_2441, signal_995}), .a ({signal_2429, signal_1059}), .c ({signal_2461, signal_1379}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1252 ( .s (signal_3301), .b ({signal_2209, signal_994}), .a ({signal_2173, signal_1058}), .c ({signal_2303, signal_1378}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1253 ( .s (signal_3301), .b ({signal_2208, signal_993}), .a ({signal_2172, signal_1057}), .c ({signal_2304, signal_1377}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1254 ( .s (signal_3301), .b ({signal_2207, signal_992}), .a ({signal_2171, signal_1056}), .c ({signal_2305, signal_1376}) ) ;
    Midori64_step2_ANF #(.low_latency(0), .pipeline(1)) cell_1255 ( .in0 ({signal_1375, signal_1374, signal_1373, signal_1372, signal_1371, signal_1370, signal_1369, signal_1368, signal_1367, signal_1366, signal_1365, signal_1364, signal_1363, signal_1362, signal_1361, signal_1360, signal_1359, signal_1358, signal_1357, signal_1356, signal_1355, signal_1354, signal_1353, signal_1352, signal_1351, signal_1350, signal_1349, signal_1348, signal_1347, signal_1346, signal_1345, signal_1344, signal_1343, signal_1342, signal_1341, signal_1340, signal_1339, signal_1338, signal_1337, signal_1336, signal_1335, signal_1334, signal_1333, signal_1332, signal_1331, signal_1330, signal_1329, signal_1328, signal_1327, signal_1326, signal_1325, signal_1324, signal_1323, signal_1322, signal_1321, signal_1320, signal_1319, signal_1318, signal_1317, signal_1316, signal_1315, signal_1314, signal_1313, signal_1312}), .in1 ({signal_1852, signal_1851, signal_1850, signal_1849, signal_1848, signal_1847, signal_1846, signal_1845, signal_1844, signal_1843, signal_1842, signal_1841, signal_1840, signal_1839, signal_1838, signal_1837, signal_1836, signal_1835, signal_1834, signal_1833, signal_1832, signal_1831, signal_1830, signal_1829, signal_1828, signal_1827, signal_1826, signal_1825, signal_1824, signal_1823, signal_1822, signal_1821, signal_1820, signal_1819, signal_1818, signal_1817, signal_1816, signal_1815, signal_1814, signal_1813, signal_1812, signal_1811, signal_1810, signal_1809, signal_1808, signal_1807, signal_1806, signal_1805, signal_1804, signal_1803, signal_1802, signal_1801, signal_1800, signal_1799, signal_1798, signal_1797, signal_1796, signal_1795, signal_1794, signal_1793, signal_1792, signal_1791, signal_1790, signal_1789}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_1311, signal_1310, signal_1309, signal_1308, signal_1307, signal_1306, signal_1305, signal_1304, signal_1303, signal_1302, signal_1301, signal_1300, signal_1299, signal_1298, signal_1297, signal_1296, signal_1295, signal_1294, signal_1293, signal_1292, signal_1291, signal_1290, signal_1289, signal_1288, signal_1287, signal_1286, signal_1285, signal_1284, signal_1283, signal_1282, signal_1281, signal_1280, signal_1279, signal_1278, signal_1277, signal_1276, signal_1275, signal_1274, signal_1273, signal_1272, signal_1271, signal_1270, signal_1269, signal_1268, signal_1267, signal_1266, signal_1265, signal_1264, signal_1263, signal_1262, signal_1261, signal_1260, signal_1259, signal_1258, signal_1257, signal_1256, signal_1255, signal_1254, signal_1253, signal_1252, signal_1251, signal_1250, signal_1249, signal_1248}), .out1 ({signal_1916, signal_1915, signal_1914, signal_1913, signal_1912, signal_1911, signal_1910, signal_1909, signal_1908, signal_1907, signal_1906, signal_1905, signal_1904, signal_1903, signal_1902, signal_1901, signal_1900, signal_1899, signal_1898, signal_1897, signal_1896, signal_1895, signal_1894, signal_1893, signal_1892, signal_1891, signal_1890, signal_1889, signal_1888, signal_1887, signal_1886, signal_1885, signal_1884, signal_1883, signal_1882, signal_1881, signal_1880, signal_1879, signal_1878, signal_1877, signal_1876, signal_1875, signal_1874, signal_1873, signal_1872, signal_1871, signal_1870, signal_1869, signal_1868, signal_1867, signal_1866, signal_1865, signal_1864, signal_1863, signal_1862, signal_1861, signal_1860, signal_1859, signal_1858, signal_1857, signal_1856, signal_1855, signal_1854, signal_1853}) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_2528), .Q (done) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_2530), .Q (signal_2531) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_2532), .Q (signal_2533) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_2534), .Q (signal_2535) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_2536), .Q (signal_2537) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_2538), .Q (signal_2539) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_2540), .Q (signal_2541) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_2542), .Q (signal_2543) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_2544), .Q (signal_2545) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_2546), .Q (signal_2547) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_2548), .Q (signal_2549) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_2550), .Q (signal_2551) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_2552), .Q (signal_2553) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_2554), .Q (signal_2555) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_2556), .Q (signal_2557) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_2558), .Q (signal_2559) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_2560), .Q (signal_2561) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_2562), .Q (signal_2563) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_2564), .Q (signal_2565) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_2566), .Q (signal_2567) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_2568), .Q (signal_2569) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_2570), .Q (signal_2571) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_2572), .Q (signal_2573) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_2574), .Q (signal_2575) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_2576), .Q (signal_2577) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_2578), .Q (signal_2579) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_2580), .Q (signal_2581) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_2582), .Q (signal_2583) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_2584), .Q (signal_2585) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_2586), .Q (signal_2587) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_2588), .Q (signal_2589) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_2590), .Q (signal_2591) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_2592), .Q (signal_2593) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_2594), .Q (signal_2595) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_2596), .Q (signal_2597) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_2598), .Q (signal_2599) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_2600), .Q (signal_2601) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_2602), .Q (signal_2603) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_2604), .Q (signal_2605) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_2606), .Q (signal_2607) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_2608), .Q (signal_2609) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_2610), .Q (signal_2611) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_2612), .Q (signal_2613) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_2614), .Q (signal_2615) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_2616), .Q (signal_2617) ) ;
    buf_clk cell_1347 ( .C (clk), .D (signal_2618), .Q (signal_2619) ) ;
    buf_clk cell_1349 ( .C (clk), .D (signal_2620), .Q (signal_2621) ) ;
    buf_clk cell_1351 ( .C (clk), .D (signal_2622), .Q (signal_2623) ) ;
    buf_clk cell_1353 ( .C (clk), .D (signal_2624), .Q (signal_2625) ) ;
    buf_clk cell_1355 ( .C (clk), .D (signal_2626), .Q (signal_2627) ) ;
    buf_clk cell_1357 ( .C (clk), .D (signal_2628), .Q (signal_2629) ) ;
    buf_clk cell_1359 ( .C (clk), .D (signal_2630), .Q (signal_2631) ) ;
    buf_clk cell_1361 ( .C (clk), .D (signal_2632), .Q (signal_2633) ) ;
    buf_clk cell_1363 ( .C (clk), .D (signal_2634), .Q (signal_2635) ) ;
    buf_clk cell_1365 ( .C (clk), .D (signal_2636), .Q (signal_2637) ) ;
    buf_clk cell_1367 ( .C (clk), .D (signal_2638), .Q (signal_2639) ) ;
    buf_clk cell_1369 ( .C (clk), .D (signal_2640), .Q (signal_2641) ) ;
    buf_clk cell_1371 ( .C (clk), .D (signal_2642), .Q (signal_2643) ) ;
    buf_clk cell_1373 ( .C (clk), .D (signal_2644), .Q (signal_2645) ) ;
    buf_clk cell_1375 ( .C (clk), .D (signal_2646), .Q (signal_2647) ) ;
    buf_clk cell_1377 ( .C (clk), .D (signal_2648), .Q (signal_2649) ) ;
    buf_clk cell_1379 ( .C (clk), .D (signal_2650), .Q (signal_2651) ) ;
    buf_clk cell_1381 ( .C (clk), .D (signal_2652), .Q (signal_2653) ) ;
    buf_clk cell_1383 ( .C (clk), .D (signal_2654), .Q (signal_2655) ) ;
    buf_clk cell_1385 ( .C (clk), .D (signal_2656), .Q (signal_2657) ) ;
    buf_clk cell_1387 ( .C (clk), .D (signal_2658), .Q (signal_2659) ) ;
    buf_clk cell_1389 ( .C (clk), .D (signal_2660), .Q (signal_2661) ) ;
    buf_clk cell_1391 ( .C (clk), .D (signal_2662), .Q (signal_2663) ) ;
    buf_clk cell_1393 ( .C (clk), .D (signal_2664), .Q (signal_2665) ) ;
    buf_clk cell_1395 ( .C (clk), .D (signal_2666), .Q (signal_2667) ) ;
    buf_clk cell_1397 ( .C (clk), .D (signal_2668), .Q (signal_2669) ) ;
    buf_clk cell_1399 ( .C (clk), .D (signal_2670), .Q (signal_2671) ) ;
    buf_clk cell_1401 ( .C (clk), .D (signal_2672), .Q (signal_2673) ) ;
    buf_clk cell_1403 ( .C (clk), .D (signal_2674), .Q (signal_2675) ) ;
    buf_clk cell_1405 ( .C (clk), .D (signal_2676), .Q (signal_2677) ) ;
    buf_clk cell_1407 ( .C (clk), .D (signal_2678), .Q (signal_2679) ) ;
    buf_clk cell_1409 ( .C (clk), .D (signal_2680), .Q (signal_2681) ) ;
    buf_clk cell_1411 ( .C (clk), .D (signal_2682), .Q (signal_2683) ) ;
    buf_clk cell_1413 ( .C (clk), .D (signal_2684), .Q (signal_2685) ) ;
    buf_clk cell_1415 ( .C (clk), .D (signal_2686), .Q (signal_2687) ) ;
    buf_clk cell_1417 ( .C (clk), .D (signal_2688), .Q (signal_2689) ) ;
    buf_clk cell_1419 ( .C (clk), .D (signal_2690), .Q (signal_2691) ) ;
    buf_clk cell_1421 ( .C (clk), .D (signal_2692), .Q (signal_2693) ) ;
    buf_clk cell_1423 ( .C (clk), .D (signal_2694), .Q (signal_2695) ) ;
    buf_clk cell_1425 ( .C (clk), .D (signal_2696), .Q (signal_2697) ) ;
    buf_clk cell_1427 ( .C (clk), .D (signal_2698), .Q (signal_2699) ) ;
    buf_clk cell_1429 ( .C (clk), .D (signal_2700), .Q (signal_2701) ) ;
    buf_clk cell_1431 ( .C (clk), .D (signal_2702), .Q (signal_2703) ) ;
    buf_clk cell_1433 ( .C (clk), .D (signal_2704), .Q (signal_2705) ) ;
    buf_clk cell_1435 ( .C (clk), .D (signal_2706), .Q (signal_2707) ) ;
    buf_clk cell_1437 ( .C (clk), .D (signal_2708), .Q (signal_2709) ) ;
    buf_clk cell_1439 ( .C (clk), .D (signal_2710), .Q (signal_2711) ) ;
    buf_clk cell_1441 ( .C (clk), .D (signal_2712), .Q (signal_2713) ) ;
    buf_clk cell_1443 ( .C (clk), .D (signal_2714), .Q (signal_2715) ) ;
    buf_clk cell_1445 ( .C (clk), .D (signal_2716), .Q (signal_2717) ) ;
    buf_clk cell_1447 ( .C (clk), .D (signal_2718), .Q (signal_2719) ) ;
    buf_clk cell_1449 ( .C (clk), .D (signal_2720), .Q (signal_2721) ) ;
    buf_clk cell_1451 ( .C (clk), .D (signal_2722), .Q (signal_2723) ) ;
    buf_clk cell_1453 ( .C (clk), .D (signal_2724), .Q (signal_2725) ) ;
    buf_clk cell_1455 ( .C (clk), .D (signal_2726), .Q (signal_2727) ) ;
    buf_clk cell_1457 ( .C (clk), .D (signal_2728), .Q (signal_2729) ) ;
    buf_clk cell_1459 ( .C (clk), .D (signal_2730), .Q (signal_2731) ) ;
    buf_clk cell_1461 ( .C (clk), .D (signal_2732), .Q (signal_2733) ) ;
    buf_clk cell_1463 ( .C (clk), .D (signal_2734), .Q (signal_2735) ) ;
    buf_clk cell_1465 ( .C (clk), .D (signal_2736), .Q (signal_2737) ) ;
    buf_clk cell_1467 ( .C (clk), .D (signal_2738), .Q (signal_2739) ) ;
    buf_clk cell_1469 ( .C (clk), .D (signal_2740), .Q (signal_2741) ) ;
    buf_clk cell_1471 ( .C (clk), .D (signal_2742), .Q (signal_2743) ) ;
    buf_clk cell_1473 ( .C (clk), .D (signal_2744), .Q (signal_2745) ) ;
    buf_clk cell_1475 ( .C (clk), .D (signal_2746), .Q (signal_2747) ) ;
    buf_clk cell_1477 ( .C (clk), .D (signal_2748), .Q (signal_2749) ) ;
    buf_clk cell_1479 ( .C (clk), .D (signal_2750), .Q (signal_2751) ) ;
    buf_clk cell_1481 ( .C (clk), .D (signal_2752), .Q (signal_2753) ) ;
    buf_clk cell_1483 ( .C (clk), .D (signal_2754), .Q (signal_2755) ) ;
    buf_clk cell_1485 ( .C (clk), .D (signal_2756), .Q (signal_2757) ) ;
    buf_clk cell_1487 ( .C (clk), .D (signal_2758), .Q (signal_2759) ) ;
    buf_clk cell_1489 ( .C (clk), .D (signal_2760), .Q (signal_2761) ) ;
    buf_clk cell_1491 ( .C (clk), .D (signal_2762), .Q (signal_2763) ) ;
    buf_clk cell_1493 ( .C (clk), .D (signal_2764), .Q (signal_2765) ) ;
    buf_clk cell_1495 ( .C (clk), .D (signal_2766), .Q (signal_2767) ) ;
    buf_clk cell_1497 ( .C (clk), .D (signal_2768), .Q (signal_2769) ) ;
    buf_clk cell_1499 ( .C (clk), .D (signal_2770), .Q (signal_2771) ) ;
    buf_clk cell_1501 ( .C (clk), .D (signal_2772), .Q (signal_2773) ) ;
    buf_clk cell_1503 ( .C (clk), .D (signal_2774), .Q (signal_2775) ) ;
    buf_clk cell_1505 ( .C (clk), .D (signal_2776), .Q (signal_2777) ) ;
    buf_clk cell_1507 ( .C (clk), .D (signal_2778), .Q (signal_2779) ) ;
    buf_clk cell_1509 ( .C (clk), .D (signal_2780), .Q (signal_2781) ) ;
    buf_clk cell_1511 ( .C (clk), .D (signal_2782), .Q (signal_2783) ) ;
    buf_clk cell_1513 ( .C (clk), .D (signal_2784), .Q (signal_2785) ) ;
    buf_clk cell_1515 ( .C (clk), .D (signal_2786), .Q (signal_2787) ) ;
    buf_clk cell_1517 ( .C (clk), .D (signal_2788), .Q (signal_2789) ) ;
    buf_clk cell_1519 ( .C (clk), .D (signal_2790), .Q (signal_2791) ) ;
    buf_clk cell_1521 ( .C (clk), .D (signal_2792), .Q (signal_2793) ) ;
    buf_clk cell_1523 ( .C (clk), .D (signal_2794), .Q (signal_2795) ) ;
    buf_clk cell_1525 ( .C (clk), .D (signal_2796), .Q (signal_2797) ) ;
    buf_clk cell_1527 ( .C (clk), .D (signal_2798), .Q (signal_2799) ) ;
    buf_clk cell_1529 ( .C (clk), .D (signal_2800), .Q (signal_2801) ) ;
    buf_clk cell_1531 ( .C (clk), .D (signal_2802), .Q (signal_2803) ) ;
    buf_clk cell_1533 ( .C (clk), .D (signal_2804), .Q (signal_2805) ) ;
    buf_clk cell_1535 ( .C (clk), .D (signal_2806), .Q (signal_2807) ) ;
    buf_clk cell_1537 ( .C (clk), .D (signal_2808), .Q (signal_2809) ) ;
    buf_clk cell_1539 ( .C (clk), .D (signal_2810), .Q (signal_2811) ) ;
    buf_clk cell_1541 ( .C (clk), .D (signal_2812), .Q (signal_2813) ) ;
    buf_clk cell_1543 ( .C (clk), .D (signal_2814), .Q (signal_2815) ) ;
    buf_clk cell_1545 ( .C (clk), .D (signal_2816), .Q (signal_2817) ) ;
    buf_clk cell_1547 ( .C (clk), .D (signal_2818), .Q (signal_2819) ) ;
    buf_clk cell_1549 ( .C (clk), .D (signal_2820), .Q (signal_2821) ) ;
    buf_clk cell_1551 ( .C (clk), .D (signal_2822), .Q (signal_2823) ) ;
    buf_clk cell_1553 ( .C (clk), .D (signal_2824), .Q (signal_2825) ) ;
    buf_clk cell_1555 ( .C (clk), .D (signal_2826), .Q (signal_2827) ) ;
    buf_clk cell_1557 ( .C (clk), .D (signal_2828), .Q (signal_2829) ) ;
    buf_clk cell_1559 ( .C (clk), .D (signal_2830), .Q (signal_2831) ) ;
    buf_clk cell_1561 ( .C (clk), .D (signal_2832), .Q (signal_2833) ) ;
    buf_clk cell_1563 ( .C (clk), .D (signal_2834), .Q (signal_2835) ) ;
    buf_clk cell_1565 ( .C (clk), .D (signal_2836), .Q (signal_2837) ) ;
    buf_clk cell_1567 ( .C (clk), .D (signal_2838), .Q (signal_2839) ) ;
    buf_clk cell_1569 ( .C (clk), .D (signal_2840), .Q (signal_2841) ) ;
    buf_clk cell_1571 ( .C (clk), .D (signal_2842), .Q (signal_2843) ) ;
    buf_clk cell_1573 ( .C (clk), .D (signal_2844), .Q (signal_2845) ) ;
    buf_clk cell_1575 ( .C (clk), .D (signal_2846), .Q (signal_2847) ) ;
    buf_clk cell_1577 ( .C (clk), .D (signal_2848), .Q (signal_2849) ) ;
    buf_clk cell_1579 ( .C (clk), .D (signal_2850), .Q (signal_2851) ) ;
    buf_clk cell_1581 ( .C (clk), .D (signal_2852), .Q (signal_2853) ) ;
    buf_clk cell_1583 ( .C (clk), .D (signal_2854), .Q (signal_2855) ) ;
    buf_clk cell_1585 ( .C (clk), .D (signal_2856), .Q (signal_2857) ) ;
    buf_clk cell_1587 ( .C (clk), .D (signal_2858), .Q (signal_2859) ) ;
    buf_clk cell_1589 ( .C (clk), .D (signal_2860), .Q (signal_2861) ) ;
    buf_clk cell_1591 ( .C (clk), .D (signal_2862), .Q (signal_2863) ) ;
    buf_clk cell_1593 ( .C (clk), .D (signal_2864), .Q (signal_2865) ) ;
    buf_clk cell_1595 ( .C (clk), .D (signal_2866), .Q (signal_2867) ) ;
    buf_clk cell_1597 ( .C (clk), .D (signal_2868), .Q (signal_2869) ) ;
    buf_clk cell_1599 ( .C (clk), .D (signal_2870), .Q (signal_2871) ) ;
    buf_clk cell_1601 ( .C (clk), .D (signal_2872), .Q (signal_2873) ) ;
    buf_clk cell_1603 ( .C (clk), .D (signal_2874), .Q (signal_2875) ) ;
    buf_clk cell_1605 ( .C (clk), .D (signal_2876), .Q (signal_2877) ) ;
    buf_clk cell_1607 ( .C (clk), .D (signal_2878), .Q (signal_2879) ) ;
    buf_clk cell_1609 ( .C (clk), .D (signal_2880), .Q (signal_2881) ) ;
    buf_clk cell_1611 ( .C (clk), .D (signal_2882), .Q (signal_2883) ) ;
    buf_clk cell_1613 ( .C (clk), .D (signal_2884), .Q (signal_2885) ) ;
    buf_clk cell_1615 ( .C (clk), .D (signal_2886), .Q (signal_2887) ) ;
    buf_clk cell_1617 ( .C (clk), .D (signal_2888), .Q (signal_2889) ) ;
    buf_clk cell_1619 ( .C (clk), .D (signal_2890), .Q (signal_2891) ) ;
    buf_clk cell_1621 ( .C (clk), .D (signal_2892), .Q (signal_2893) ) ;
    buf_clk cell_1623 ( .C (clk), .D (signal_2894), .Q (signal_2895) ) ;
    buf_clk cell_1625 ( .C (clk), .D (signal_2896), .Q (signal_2897) ) ;
    buf_clk cell_1627 ( .C (clk), .D (signal_2898), .Q (signal_2899) ) ;
    buf_clk cell_1629 ( .C (clk), .D (signal_2900), .Q (signal_2901) ) ;
    buf_clk cell_1631 ( .C (clk), .D (signal_2902), .Q (signal_2903) ) ;
    buf_clk cell_1633 ( .C (clk), .D (signal_2904), .Q (signal_2905) ) ;
    buf_clk cell_1635 ( .C (clk), .D (signal_2906), .Q (signal_2907) ) ;
    buf_clk cell_1637 ( .C (clk), .D (signal_2908), .Q (signal_2909) ) ;
    buf_clk cell_1639 ( .C (clk), .D (signal_2910), .Q (signal_2911) ) ;
    buf_clk cell_1641 ( .C (clk), .D (signal_2912), .Q (signal_2913) ) ;
    buf_clk cell_1643 ( .C (clk), .D (signal_2914), .Q (signal_2915) ) ;
    buf_clk cell_1645 ( .C (clk), .D (signal_2916), .Q (signal_2917) ) ;
    buf_clk cell_1647 ( .C (clk), .D (signal_2918), .Q (signal_2919) ) ;
    buf_clk cell_1649 ( .C (clk), .D (signal_2920), .Q (signal_2921) ) ;
    buf_clk cell_1651 ( .C (clk), .D (signal_2922), .Q (signal_2923) ) ;
    buf_clk cell_1653 ( .C (clk), .D (signal_2924), .Q (signal_2925) ) ;
    buf_clk cell_1655 ( .C (clk), .D (signal_2926), .Q (signal_2927) ) ;
    buf_clk cell_1657 ( .C (clk), .D (signal_2928), .Q (signal_2929) ) ;
    buf_clk cell_1659 ( .C (clk), .D (signal_2930), .Q (signal_2931) ) ;
    buf_clk cell_1661 ( .C (clk), .D (signal_2932), .Q (signal_2933) ) ;
    buf_clk cell_1663 ( .C (clk), .D (signal_2934), .Q (signal_2935) ) ;
    buf_clk cell_1665 ( .C (clk), .D (signal_2936), .Q (signal_2937) ) ;
    buf_clk cell_1667 ( .C (clk), .D (signal_2938), .Q (signal_2939) ) ;
    buf_clk cell_1669 ( .C (clk), .D (signal_2940), .Q (signal_2941) ) ;
    buf_clk cell_1671 ( .C (clk), .D (signal_2942), .Q (signal_2943) ) ;
    buf_clk cell_1673 ( .C (clk), .D (signal_2944), .Q (signal_2945) ) ;
    buf_clk cell_1675 ( .C (clk), .D (signal_2946), .Q (signal_2947) ) ;
    buf_clk cell_1677 ( .C (clk), .D (signal_2948), .Q (signal_2949) ) ;
    buf_clk cell_1679 ( .C (clk), .D (signal_2950), .Q (signal_2951) ) ;
    buf_clk cell_1681 ( .C (clk), .D (signal_2952), .Q (signal_2953) ) ;
    buf_clk cell_1683 ( .C (clk), .D (signal_2954), .Q (signal_2955) ) ;
    buf_clk cell_1685 ( .C (clk), .D (signal_2956), .Q (signal_2957) ) ;
    buf_clk cell_1687 ( .C (clk), .D (signal_2958), .Q (signal_2959) ) ;
    buf_clk cell_1689 ( .C (clk), .D (signal_2960), .Q (signal_2961) ) ;
    buf_clk cell_1691 ( .C (clk), .D (signal_2962), .Q (signal_2963) ) ;
    buf_clk cell_1693 ( .C (clk), .D (signal_2964), .Q (signal_2965) ) ;
    buf_clk cell_1695 ( .C (clk), .D (signal_2966), .Q (signal_2967) ) ;
    buf_clk cell_1697 ( .C (clk), .D (signal_2968), .Q (signal_2969) ) ;
    buf_clk cell_1699 ( .C (clk), .D (signal_2970), .Q (signal_2971) ) ;
    buf_clk cell_1701 ( .C (clk), .D (signal_2972), .Q (signal_2973) ) ;
    buf_clk cell_1703 ( .C (clk), .D (signal_2974), .Q (signal_2975) ) ;
    buf_clk cell_1705 ( .C (clk), .D (signal_2976), .Q (signal_2977) ) ;
    buf_clk cell_1707 ( .C (clk), .D (signal_2978), .Q (signal_2979) ) ;
    buf_clk cell_1709 ( .C (clk), .D (signal_2980), .Q (signal_2981) ) ;
    buf_clk cell_1711 ( .C (clk), .D (signal_2982), .Q (signal_2983) ) ;
    buf_clk cell_1713 ( .C (clk), .D (signal_2984), .Q (signal_2985) ) ;
    buf_clk cell_1715 ( .C (clk), .D (signal_2986), .Q (signal_2987) ) ;
    buf_clk cell_1717 ( .C (clk), .D (signal_2988), .Q (signal_2989) ) ;
    buf_clk cell_1719 ( .C (clk), .D (signal_2990), .Q (signal_2991) ) ;
    buf_clk cell_1721 ( .C (clk), .D (signal_2992), .Q (signal_2993) ) ;
    buf_clk cell_1723 ( .C (clk), .D (signal_2994), .Q (signal_2995) ) ;
    buf_clk cell_1725 ( .C (clk), .D (signal_2996), .Q (signal_2997) ) ;
    buf_clk cell_1727 ( .C (clk), .D (signal_2998), .Q (signal_2999) ) ;
    buf_clk cell_1729 ( .C (clk), .D (signal_3000), .Q (signal_3001) ) ;
    buf_clk cell_1731 ( .C (clk), .D (signal_3002), .Q (signal_3003) ) ;
    buf_clk cell_1733 ( .C (clk), .D (signal_3004), .Q (signal_3005) ) ;
    buf_clk cell_1735 ( .C (clk), .D (signal_3006), .Q (signal_3007) ) ;
    buf_clk cell_1737 ( .C (clk), .D (signal_3008), .Q (signal_3009) ) ;
    buf_clk cell_1739 ( .C (clk), .D (signal_3010), .Q (signal_3011) ) ;
    buf_clk cell_1741 ( .C (clk), .D (signal_3012), .Q (signal_3013) ) ;
    buf_clk cell_1743 ( .C (clk), .D (signal_3014), .Q (signal_3015) ) ;
    buf_clk cell_1745 ( .C (clk), .D (signal_3016), .Q (signal_3017) ) ;
    buf_clk cell_1747 ( .C (clk), .D (signal_3018), .Q (signal_3019) ) ;
    buf_clk cell_1749 ( .C (clk), .D (signal_3020), .Q (signal_3021) ) ;
    buf_clk cell_1751 ( .C (clk), .D (signal_3022), .Q (signal_3023) ) ;
    buf_clk cell_1753 ( .C (clk), .D (signal_3024), .Q (signal_3025) ) ;
    buf_clk cell_1755 ( .C (clk), .D (signal_3026), .Q (signal_3027) ) ;
    buf_clk cell_1757 ( .C (clk), .D (signal_3028), .Q (signal_3029) ) ;
    buf_clk cell_1759 ( .C (clk), .D (signal_3030), .Q (signal_3031) ) ;
    buf_clk cell_1761 ( .C (clk), .D (signal_3032), .Q (signal_3033) ) ;
    buf_clk cell_1763 ( .C (clk), .D (signal_3034), .Q (signal_3035) ) ;
    buf_clk cell_1765 ( .C (clk), .D (signal_3036), .Q (signal_3037) ) ;
    buf_clk cell_1767 ( .C (clk), .D (signal_3038), .Q (signal_3039) ) ;
    buf_clk cell_1769 ( .C (clk), .D (signal_3040), .Q (signal_3041) ) ;
    buf_clk cell_1771 ( .C (clk), .D (signal_3042), .Q (signal_3043) ) ;
    buf_clk cell_1773 ( .C (clk), .D (signal_3044), .Q (signal_3045) ) ;
    buf_clk cell_1775 ( .C (clk), .D (signal_3046), .Q (signal_3047) ) ;
    buf_clk cell_1777 ( .C (clk), .D (signal_3048), .Q (signal_3049) ) ;
    buf_clk cell_1779 ( .C (clk), .D (signal_3050), .Q (signal_3051) ) ;
    buf_clk cell_1781 ( .C (clk), .D (signal_3052), .Q (signal_3053) ) ;
    buf_clk cell_1783 ( .C (clk), .D (signal_3054), .Q (signal_3055) ) ;
    buf_clk cell_1785 ( .C (clk), .D (signal_3056), .Q (signal_3057) ) ;
    buf_clk cell_1787 ( .C (clk), .D (signal_3058), .Q (signal_3059) ) ;
    buf_clk cell_1789 ( .C (clk), .D (signal_3060), .Q (signal_3061) ) ;
    buf_clk cell_1791 ( .C (clk), .D (signal_3062), .Q (signal_3063) ) ;
    buf_clk cell_1793 ( .C (clk), .D (signal_3064), .Q (signal_3065) ) ;
    buf_clk cell_1795 ( .C (clk), .D (signal_3066), .Q (signal_3067) ) ;
    buf_clk cell_1797 ( .C (clk), .D (signal_3068), .Q (signal_3069) ) ;
    buf_clk cell_1799 ( .C (clk), .D (signal_3070), .Q (signal_3071) ) ;
    buf_clk cell_1801 ( .C (clk), .D (signal_3072), .Q (signal_3073) ) ;
    buf_clk cell_1803 ( .C (clk), .D (signal_3074), .Q (signal_3075) ) ;
    buf_clk cell_1805 ( .C (clk), .D (signal_3076), .Q (signal_3077) ) ;
    buf_clk cell_1807 ( .C (clk), .D (signal_3078), .Q (signal_3079) ) ;
    buf_clk cell_1809 ( .C (clk), .D (signal_3080), .Q (signal_3081) ) ;
    buf_clk cell_1811 ( .C (clk), .D (signal_3082), .Q (signal_3083) ) ;
    buf_clk cell_1813 ( .C (clk), .D (signal_3084), .Q (signal_3085) ) ;
    buf_clk cell_1815 ( .C (clk), .D (signal_3086), .Q (signal_3087) ) ;
    buf_clk cell_1817 ( .C (clk), .D (signal_3088), .Q (signal_3089) ) ;
    buf_clk cell_1819 ( .C (clk), .D (signal_3090), .Q (signal_3091) ) ;
    buf_clk cell_1821 ( .C (clk), .D (signal_3092), .Q (signal_3093) ) ;
    buf_clk cell_1823 ( .C (clk), .D (signal_3094), .Q (signal_3095) ) ;
    buf_clk cell_1825 ( .C (clk), .D (signal_3096), .Q (signal_3097) ) ;
    buf_clk cell_1827 ( .C (clk), .D (signal_3098), .Q (signal_3099) ) ;
    buf_clk cell_1829 ( .C (clk), .D (signal_3100), .Q (signal_3101) ) ;
    buf_clk cell_1831 ( .C (clk), .D (signal_3102), .Q (signal_3103) ) ;
    buf_clk cell_1833 ( .C (clk), .D (signal_3104), .Q (signal_3105) ) ;
    buf_clk cell_1835 ( .C (clk), .D (signal_3106), .Q (signal_3107) ) ;
    buf_clk cell_1837 ( .C (clk), .D (signal_3108), .Q (signal_3109) ) ;
    buf_clk cell_1839 ( .C (clk), .D (signal_3110), .Q (signal_3111) ) ;
    buf_clk cell_1841 ( .C (clk), .D (signal_3112), .Q (signal_3113) ) ;
    buf_clk cell_1843 ( .C (clk), .D (signal_3114), .Q (signal_3115) ) ;
    buf_clk cell_1845 ( .C (clk), .D (signal_3116), .Q (signal_3117) ) ;
    buf_clk cell_1847 ( .C (clk), .D (signal_3118), .Q (signal_3119) ) ;
    buf_clk cell_1849 ( .C (clk), .D (signal_3120), .Q (signal_3121) ) ;
    buf_clk cell_1851 ( .C (clk), .D (signal_3122), .Q (signal_3123) ) ;
    buf_clk cell_1853 ( .C (clk), .D (signal_3124), .Q (signal_3125) ) ;
    buf_clk cell_1855 ( .C (clk), .D (signal_3126), .Q (signal_3127) ) ;
    buf_clk cell_1857 ( .C (clk), .D (signal_3128), .Q (signal_3129) ) ;
    buf_clk cell_1859 ( .C (clk), .D (signal_3130), .Q (signal_3131) ) ;
    buf_clk cell_1861 ( .C (clk), .D (signal_3132), .Q (signal_3133) ) ;
    buf_clk cell_1863 ( .C (clk), .D (signal_3134), .Q (signal_3135) ) ;
    buf_clk cell_1865 ( .C (clk), .D (signal_3136), .Q (signal_3137) ) ;
    buf_clk cell_1867 ( .C (clk), .D (signal_3138), .Q (signal_3139) ) ;
    buf_clk cell_1869 ( .C (clk), .D (signal_3140), .Q (signal_3141) ) ;
    buf_clk cell_1871 ( .C (clk), .D (signal_3142), .Q (signal_3143) ) ;
    buf_clk cell_1873 ( .C (clk), .D (signal_3144), .Q (signal_3145) ) ;
    buf_clk cell_1875 ( .C (clk), .D (signal_3146), .Q (signal_3147) ) ;
    buf_clk cell_1877 ( .C (clk), .D (signal_3148), .Q (signal_3149) ) ;
    buf_clk cell_1879 ( .C (clk), .D (signal_3150), .Q (signal_3151) ) ;
    buf_clk cell_1881 ( .C (clk), .D (signal_3152), .Q (signal_3153) ) ;
    buf_clk cell_1883 ( .C (clk), .D (signal_3154), .Q (signal_3155) ) ;
    buf_clk cell_1885 ( .C (clk), .D (signal_3156), .Q (signal_3157) ) ;
    buf_clk cell_1887 ( .C (clk), .D (signal_3158), .Q (signal_3159) ) ;
    buf_clk cell_1889 ( .C (clk), .D (signal_3160), .Q (signal_3161) ) ;
    buf_clk cell_1891 ( .C (clk), .D (signal_3162), .Q (signal_3163) ) ;
    buf_clk cell_1893 ( .C (clk), .D (signal_3164), .Q (signal_3165) ) ;
    buf_clk cell_1895 ( .C (clk), .D (signal_3166), .Q (signal_3167) ) ;
    buf_clk cell_1897 ( .C (clk), .D (signal_3168), .Q (signal_3169) ) ;
    buf_clk cell_1899 ( .C (clk), .D (signal_3170), .Q (signal_3171) ) ;
    buf_clk cell_1901 ( .C (clk), .D (signal_3172), .Q (signal_3173) ) ;
    buf_clk cell_1903 ( .C (clk), .D (signal_3174), .Q (signal_3175) ) ;
    buf_clk cell_1905 ( .C (clk), .D (signal_3176), .Q (signal_3177) ) ;
    buf_clk cell_1907 ( .C (clk), .D (signal_3178), .Q (signal_3179) ) ;
    buf_clk cell_1909 ( .C (clk), .D (signal_3180), .Q (signal_3181) ) ;
    buf_clk cell_1911 ( .C (clk), .D (signal_3182), .Q (signal_3183) ) ;
    buf_clk cell_1913 ( .C (clk), .D (signal_3184), .Q (signal_3185) ) ;
    buf_clk cell_1915 ( .C (clk), .D (signal_3186), .Q (signal_3187) ) ;
    buf_clk cell_1917 ( .C (clk), .D (signal_3188), .Q (signal_3189) ) ;
    buf_clk cell_1919 ( .C (clk), .D (signal_3190), .Q (signal_3191) ) ;
    buf_clk cell_1921 ( .C (clk), .D (signal_3192), .Q (signal_3193) ) ;
    buf_clk cell_1923 ( .C (clk), .D (signal_3194), .Q (signal_3195) ) ;
    buf_clk cell_1925 ( .C (clk), .D (signal_3196), .Q (signal_3197) ) ;
    buf_clk cell_1927 ( .C (clk), .D (signal_3198), .Q (signal_3199) ) ;
    buf_clk cell_1929 ( .C (clk), .D (signal_3200), .Q (signal_3201) ) ;
    buf_clk cell_1931 ( .C (clk), .D (signal_3202), .Q (signal_3203) ) ;
    buf_clk cell_1933 ( .C (clk), .D (signal_3204), .Q (signal_3205) ) ;
    buf_clk cell_1935 ( .C (clk), .D (signal_3206), .Q (signal_3207) ) ;
    buf_clk cell_1937 ( .C (clk), .D (signal_3208), .Q (signal_3209) ) ;
    buf_clk cell_1939 ( .C (clk), .D (signal_3210), .Q (signal_3211) ) ;
    buf_clk cell_1941 ( .C (clk), .D (signal_3212), .Q (signal_3213) ) ;
    buf_clk cell_1943 ( .C (clk), .D (signal_3214), .Q (signal_3215) ) ;
    buf_clk cell_1945 ( .C (clk), .D (signal_3216), .Q (signal_3217) ) ;
    buf_clk cell_1947 ( .C (clk), .D (signal_3218), .Q (signal_3219) ) ;
    buf_clk cell_1949 ( .C (clk), .D (signal_3220), .Q (signal_3221) ) ;
    buf_clk cell_1951 ( .C (clk), .D (signal_3222), .Q (signal_3223) ) ;
    buf_clk cell_1953 ( .C (clk), .D (signal_3224), .Q (signal_3225) ) ;
    buf_clk cell_1955 ( .C (clk), .D (signal_3226), .Q (signal_3227) ) ;
    buf_clk cell_1957 ( .C (clk), .D (signal_3228), .Q (signal_3229) ) ;
    buf_clk cell_1959 ( .C (clk), .D (signal_3230), .Q (signal_3231) ) ;
    buf_clk cell_1961 ( .C (clk), .D (signal_3232), .Q (signal_3233) ) ;
    buf_clk cell_1963 ( .C (clk), .D (signal_3234), .Q (signal_3235) ) ;
    buf_clk cell_1965 ( .C (clk), .D (signal_3236), .Q (signal_3237) ) ;
    buf_clk cell_1967 ( .C (clk), .D (signal_3238), .Q (signal_3239) ) ;
    buf_clk cell_1969 ( .C (clk), .D (signal_3240), .Q (signal_3241) ) ;
    buf_clk cell_1971 ( .C (clk), .D (signal_3242), .Q (signal_3243) ) ;
    buf_clk cell_1973 ( .C (clk), .D (signal_3244), .Q (signal_3245) ) ;
    buf_clk cell_1975 ( .C (clk), .D (signal_3246), .Q (signal_3247) ) ;
    buf_clk cell_1977 ( .C (clk), .D (signal_3248), .Q (signal_3249) ) ;
    buf_clk cell_1979 ( .C (clk), .D (signal_3250), .Q (signal_3251) ) ;
    buf_clk cell_1981 ( .C (clk), .D (signal_3252), .Q (signal_3253) ) ;
    buf_clk cell_1983 ( .C (clk), .D (signal_3254), .Q (signal_3255) ) ;
    buf_clk cell_1985 ( .C (clk), .D (signal_3256), .Q (signal_3257) ) ;
    buf_clk cell_1987 ( .C (clk), .D (signal_3258), .Q (signal_3259) ) ;
    buf_clk cell_1989 ( .C (clk), .D (signal_3260), .Q (signal_3261) ) ;
    buf_clk cell_1991 ( .C (clk), .D (signal_3262), .Q (signal_3263) ) ;
    buf_clk cell_1993 ( .C (clk), .D (signal_3264), .Q (signal_3265) ) ;
    buf_clk cell_1995 ( .C (clk), .D (signal_3266), .Q (signal_3267) ) ;
    buf_clk cell_1997 ( .C (clk), .D (signal_3268), .Q (signal_3269) ) ;
    buf_clk cell_1999 ( .C (clk), .D (signal_3270), .Q (signal_3271) ) ;
    buf_clk cell_2001 ( .C (clk), .D (signal_3272), .Q (signal_3273) ) ;
    buf_clk cell_2003 ( .C (clk), .D (signal_3274), .Q (signal_3275) ) ;
    buf_clk cell_2005 ( .C (clk), .D (signal_3276), .Q (signal_3277) ) ;
    buf_clk cell_2007 ( .C (clk), .D (signal_3278), .Q (signal_3279) ) ;
    buf_clk cell_2009 ( .C (clk), .D (signal_3280), .Q (signal_3281) ) ;
    buf_clk cell_2011 ( .C (clk), .D (signal_3282), .Q (signal_3283) ) ;
    buf_clk cell_2013 ( .C (clk), .D (signal_3284), .Q (signal_3285) ) ;
    buf_clk cell_2015 ( .C (clk), .D (signal_3286), .Q (signal_3287) ) ;
    buf_clk cell_2017 ( .C (clk), .D (signal_3288), .Q (signal_3289) ) ;
    buf_clk cell_2019 ( .C (clk), .D (signal_3290), .Q (signal_3291) ) ;
    buf_clk cell_2021 ( .C (clk), .D (signal_3292), .Q (signal_3293) ) ;
    buf_clk cell_2023 ( .C (clk), .D (signal_3294), .Q (signal_3295) ) ;
    buf_clk cell_2025 ( .C (clk), .D (signal_3296), .Q (signal_3297) ) ;
    buf_clk cell_2027 ( .C (clk), .D (signal_3298), .Q (signal_3299) ) ;
    buf_clk cell_2029 ( .C (clk), .D (signal_3300), .Q (signal_3301) ) ;
    buf_clk cell_2031 ( .C (clk), .D (signal_3302), .Q (signal_3303) ) ;
    buf_clk cell_2033 ( .C (clk), .D (signal_3304), .Q (signal_3305) ) ;
    buf_clk cell_2035 ( .C (clk), .D (signal_3306), .Q (signal_3307) ) ;
    buf_clk cell_2037 ( .C (clk), .D (signal_3308), .Q (signal_3309) ) ;

    /* register cells */
    DFF_X1 cell_82 ( .CK (clk), .D (signal_3303), .Q (signal_927), .QN () ) ;
    DFF_X1 cell_84 ( .CK (clk), .D (signal_3305), .Q (signal_926), .QN () ) ;
    DFF_X1 cell_86 ( .CK (clk), .D (signal_3307), .Q (signal_925), .QN () ) ;
    DFF_X1 cell_88 ( .CK (clk), .D (signal_3309), .Q (signal_924), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_537 ( .clk (clk), .D ({signal_2443, signal_460}), .Q ({signal_1852, signal_1375}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_540 ( .clk (clk), .D ({signal_2258, signal_462}), .Q ({signal_1851, signal_1374}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_543 ( .clk (clk), .D ({signal_2259, signal_464}), .Q ({signal_1850, signal_1373}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_546 ( .clk (clk), .D ({signal_2260, signal_466}), .Q ({signal_1849, signal_1372}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_549 ( .clk (clk), .D ({signal_2444, signal_468}), .Q ({signal_1848, signal_1371}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_552 ( .clk (clk), .D ({signal_2261, signal_470}), .Q ({signal_1847, signal_1370}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_555 ( .clk (clk), .D ({signal_2262, signal_472}), .Q ({signal_1846, signal_1369}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_558 ( .clk (clk), .D ({signal_2263, signal_474}), .Q ({signal_1845, signal_1368}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_561 ( .clk (clk), .D ({signal_2445, signal_476}), .Q ({signal_1844, signal_1367}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_564 ( .clk (clk), .D ({signal_2320, signal_478}), .Q ({signal_1843, signal_1366}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_567 ( .clk (clk), .D ({signal_2321, signal_480}), .Q ({signal_1842, signal_1365}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_570 ( .clk (clk), .D ({signal_2322, signal_482}), .Q ({signal_1841, signal_1364}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_573 ( .clk (clk), .D ({signal_2446, signal_484}), .Q ({signal_1840, signal_1363}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_576 ( .clk (clk), .D ({signal_2323, signal_486}), .Q ({signal_1839, signal_1362}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_579 ( .clk (clk), .D ({signal_2324, signal_488}), .Q ({signal_1838, signal_1361}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_582 ( .clk (clk), .D ({signal_2325, signal_490}), .Q ({signal_1837, signal_1360}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_585 ( .clk (clk), .D ({signal_2457, signal_492}), .Q ({signal_1836, signal_1359}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_588 ( .clk (clk), .D ({signal_2326, signal_494}), .Q ({signal_1835, signal_1358}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_591 ( .clk (clk), .D ({signal_2327, signal_496}), .Q ({signal_1834, signal_1357}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_594 ( .clk (clk), .D ({signal_2328, signal_498}), .Q ({signal_1833, signal_1356}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_597 ( .clk (clk), .D ({signal_2458, signal_500}), .Q ({signal_1832, signal_1355}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_600 ( .clk (clk), .D ({signal_2329, signal_502}), .Q ({signal_1831, signal_1354}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_603 ( .clk (clk), .D ({signal_2330, signal_504}), .Q ({signal_1830, signal_1353}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_606 ( .clk (clk), .D ({signal_2331, signal_506}), .Q ({signal_1829, signal_1352}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_609 ( .clk (clk), .D ({signal_2447, signal_508}), .Q ({signal_1828, signal_1351}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_612 ( .clk (clk), .D ({signal_2332, signal_510}), .Q ({signal_1827, signal_1350}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_615 ( .clk (clk), .D ({signal_2333, signal_512}), .Q ({signal_1826, signal_1349}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_618 ( .clk (clk), .D ({signal_2334, signal_514}), .Q ({signal_1825, signal_1348}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_621 ( .clk (clk), .D ({signal_2448, signal_516}), .Q ({signal_1824, signal_1347}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_624 ( .clk (clk), .D ({signal_2335, signal_518}), .Q ({signal_1823, signal_1346}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_627 ( .clk (clk), .D ({signal_2336, signal_520}), .Q ({signal_1822, signal_1345}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_630 ( .clk (clk), .D ({signal_2337, signal_522}), .Q ({signal_1821, signal_1344}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_633 ( .clk (clk), .D ({signal_2449, signal_524}), .Q ({signal_1820, signal_1343}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_636 ( .clk (clk), .D ({signal_2338, signal_526}), .Q ({signal_1819, signal_1342}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_639 ( .clk (clk), .D ({signal_2339, signal_528}), .Q ({signal_1818, signal_1341}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_642 ( .clk (clk), .D ({signal_2340, signal_530}), .Q ({signal_1817, signal_1340}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_645 ( .clk (clk), .D ({signal_2450, signal_532}), .Q ({signal_1816, signal_1339}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_648 ( .clk (clk), .D ({signal_2341, signal_534}), .Q ({signal_1815, signal_1338}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_651 ( .clk (clk), .D ({signal_2342, signal_536}), .Q ({signal_1814, signal_1337}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_654 ( .clk (clk), .D ({signal_2343, signal_538}), .Q ({signal_1813, signal_1336}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_657 ( .clk (clk), .D ({signal_2451, signal_540}), .Q ({signal_1812, signal_1335}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_660 ( .clk (clk), .D ({signal_2344, signal_542}), .Q ({signal_1811, signal_1334}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_663 ( .clk (clk), .D ({signal_2345, signal_544}), .Q ({signal_1810, signal_1333}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_666 ( .clk (clk), .D ({signal_2346, signal_546}), .Q ({signal_1809, signal_1332}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_669 ( .clk (clk), .D ({signal_2452, signal_548}), .Q ({signal_1808, signal_1331}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_672 ( .clk (clk), .D ({signal_2347, signal_550}), .Q ({signal_1807, signal_1330}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_675 ( .clk (clk), .D ({signal_2348, signal_552}), .Q ({signal_1806, signal_1329}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_678 ( .clk (clk), .D ({signal_2349, signal_554}), .Q ({signal_1805, signal_1328}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_681 ( .clk (clk), .D ({signal_2453, signal_556}), .Q ({signal_1804, signal_1327}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_684 ( .clk (clk), .D ({signal_2350, signal_558}), .Q ({signal_1803, signal_1326}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_687 ( .clk (clk), .D ({signal_2351, signal_560}), .Q ({signal_1802, signal_1325}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_690 ( .clk (clk), .D ({signal_2352, signal_562}), .Q ({signal_1801, signal_1324}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_693 ( .clk (clk), .D ({signal_2459, signal_564}), .Q ({signal_1800, signal_1323}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_696 ( .clk (clk), .D ({signal_2353, signal_566}), .Q ({signal_1799, signal_1322}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_699 ( .clk (clk), .D ({signal_2354, signal_568}), .Q ({signal_1798, signal_1321}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_702 ( .clk (clk), .D ({signal_2355, signal_570}), .Q ({signal_1797, signal_1320}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_705 ( .clk (clk), .D ({signal_2462, signal_572}), .Q ({signal_1796, signal_1319}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_708 ( .clk (clk), .D ({signal_2356, signal_574}), .Q ({signal_1795, signal_1318}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_711 ( .clk (clk), .D ({signal_2357, signal_576}), .Q ({signal_1794, signal_1317}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_714 ( .clk (clk), .D ({signal_2358, signal_578}), .Q ({signal_1793, signal_1316}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_717 ( .clk (clk), .D ({signal_2463, signal_580}), .Q ({signal_1792, signal_1315}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_720 ( .clk (clk), .D ({signal_2359, signal_582}), .Q ({signal_1791, signal_1314}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_723 ( .clk (clk), .D ({signal_2360, signal_584}), .Q ({signal_1790, signal_1313}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_726 ( .clk (clk), .D ({signal_2361, signal_586}), .Q ({signal_1789, signal_1312}) ) ;
endmodule
