/* modified netlist. Source: module sbox in file Designs/AESSbox/Canright/AGEMA/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_GHPCLL_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [159:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire sbe_n10 ;
    wire sbe_n9 ;
    wire sbe_n8 ;
    wire sbe_n7 ;
    wire sbe_n6 ;
    wire sbe_n5 ;
    wire sbe_n4 ;
    wire sbe_n3 ;
    wire sbe_n12 ;
    wire sbe_n11 ;
    wire sbe_n2 ;
    wire sbe_n1 ;
    wire sbe_n25 ;
    wire sbe_n24 ;
    wire sbe_n23 ;
    wire sbe_n22 ;
    wire sbe_n21 ;
    wire sbe_n20 ;
    wire sbe_n19 ;
    wire sbe_n18 ;
    wire sbe_n17 ;
    wire sbe_n16 ;
    wire sbe_n15 ;
    wire sbe_n14 ;
    wire sbe_D_0_ ;
    wire sbe_D_2_ ;
    wire sbe_D_3_ ;
    wire sbe_D_5_ ;
    wire sbe_D_6_ ;
    wire sbe_C_0_ ;
    wire sbe_C_1_ ;
    wire sbe_C_2_ ;
    wire sbe_C_3_ ;
    wire sbe_C_4_ ;
    wire sbe_C_5_ ;
    wire sbe_C_6_ ;
    wire sbe_C_7_ ;
    wire sbe_Y_0_ ;
    wire sbe_Y_1_ ;
    wire sbe_Y_2_ ;
    wire sbe_Y_4_ ;
    wire sbe_Y_5_ ;
    wire sbe_Y_6_ ;
    wire sbe_B_3_ ;
    wire sbe_B_6_ ;
    wire sbe_sel_in_m7_n8 ;
    wire sbe_sel_in_m6_n8 ;
    wire sbe_sel_in_m5_n8 ;
    wire sbe_sel_in_m4_n8 ;
    wire sbe_sel_in_m3_n8 ;
    wire sbe_sel_in_m2_n8 ;
    wire sbe_sel_in_m1_n8 ;
    wire sbe_sel_in_m0_n8 ;
    wire sbe_inv_n21 ;
    wire sbe_inv_n20 ;
    wire sbe_inv_n19 ;
    wire sbe_inv_n18 ;
    wire sbe_inv_n17 ;
    wire sbe_inv_n16 ;
    wire sbe_inv_n15 ;
    wire sbe_inv_n14 ;
    wire sbe_inv_n13 ;
    wire sbe_inv_n12 ;
    wire sbe_inv_n11 ;
    wire sbe_inv_n10 ;
    wire sbe_inv_n9 ;
    wire sbe_inv_n8 ;
    wire sbe_inv_n7 ;
    wire sbe_inv_n6 ;
    wire sbe_inv_n5 ;
    wire sbe_inv_n4 ;
    wire sbe_inv_n3 ;
    wire sbe_inv_n2 ;
    wire sbe_inv_dd ;
    wire sbe_inv_dh ;
    wire sbe_inv_dl ;
    wire sbe_inv_sd_0_ ;
    wire sbe_inv_sd_1_ ;
    wire sbe_inv_d_0_ ;
    wire sbe_inv_d_1_ ;
    wire sbe_inv_d_2_ ;
    wire sbe_inv_d_3_ ;
    wire sbe_inv_bb ;
    wire sbe_inv_bh ;
    wire sbe_inv_bl ;
    wire sbe_inv_aa ;
    wire sbe_inv_ah ;
    wire sbe_inv_al ;
    wire sbe_inv_sb_0_ ;
    wire sbe_inv_sb_1_ ;
    wire sbe_inv_sa_0_ ;
    wire sbe_inv_sa_1_ ;
    wire sbe_inv_dinv_n4 ;
    wire sbe_inv_dinv_n3 ;
    wire sbe_inv_dinv_n2 ;
    wire sbe_inv_dinv_n1 ;
    wire sbe_inv_dinv_sd ;
    wire sbe_inv_dinv_d_0_ ;
    wire sbe_inv_dinv_d_1_ ;
    wire sbe_inv_dinv_sb ;
    wire sbe_inv_dinv_sa ;
    wire sbe_inv_dinv_pmul_n9 ;
    wire sbe_inv_dinv_pmul_n8 ;
    wire sbe_inv_dinv_pmul_n7 ;
    wire sbe_inv_dinv_qmul_n9 ;
    wire sbe_inv_dinv_qmul_n8 ;
    wire sbe_inv_dinv_qmul_n7 ;
    wire sbe_inv_pmul_p_0_ ;
    wire sbe_inv_pmul_p_1_ ;
    wire sbe_inv_pmul_himul_n9 ;
    wire sbe_inv_pmul_himul_n8 ;
    wire sbe_inv_pmul_himul_n7 ;
    wire sbe_inv_pmul_lomul_n9 ;
    wire sbe_inv_pmul_lomul_n8 ;
    wire sbe_inv_pmul_lomul_n7 ;
    wire sbe_inv_pmul_summul_n9 ;
    wire sbe_inv_pmul_summul_n8 ;
    wire sbe_inv_pmul_summul_n7 ;
    wire sbe_inv_qmul_p_0_ ;
    wire sbe_inv_qmul_p_1_ ;
    wire sbe_inv_qmul_himul_n9 ;
    wire sbe_inv_qmul_himul_n8 ;
    wire sbe_inv_qmul_himul_n7 ;
    wire sbe_inv_qmul_lomul_n9 ;
    wire sbe_inv_qmul_lomul_n8 ;
    wire sbe_inv_qmul_lomul_n7 ;
    wire sbe_inv_qmul_summul_n9 ;
    wire sbe_inv_qmul_summul_n8 ;
    wire sbe_inv_qmul_summul_n7 ;
    wire sbe_sel_out_m7_n8 ;
    wire sbe_sel_out_m6_n8 ;
    wire sbe_sel_out_m5_n8 ;
    wire sbe_sel_out_m4_n8 ;
    wire sbe_sel_out_m3_n8 ;
    wire sbe_sel_out_m2_n8 ;
    wire sbe_sel_out_m1_n8 ;
    wire sbe_sel_out_m0_n8 ;
    wire [7:0] O ;
    wire [6:3] sbe_X ;
    wire [7:0] sbe_Z ;
    wire [3:0] sbe_inv_c ;
    wire [1:0] sbe_inv_pmul_pl ;
    wire [1:0] sbe_inv_pmul_ph ;
    wire [1:0] sbe_inv_qmul_pl ;
    wire [1:0] sbe_inv_qmul_ph ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;
    wire new_AGEMA_signal_593 ;
    wire new_AGEMA_signal_594 ;
    wire new_AGEMA_signal_595 ;
    wire new_AGEMA_signal_596 ;
    wire new_AGEMA_signal_597 ;
    wire new_AGEMA_signal_598 ;
    wire new_AGEMA_signal_599 ;
    wire new_AGEMA_signal_600 ;
    wire new_AGEMA_signal_601 ;
    wire new_AGEMA_signal_602 ;
    wire new_AGEMA_signal_603 ;
    wire new_AGEMA_signal_604 ;
    wire new_AGEMA_signal_605 ;
    wire new_AGEMA_signal_606 ;
    wire new_AGEMA_signal_607 ;
    wire new_AGEMA_signal_608 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;

    /* cells in depth 0 */
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U39 ( .a ({X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_211, sbe_n25}), .c ({new_AGEMA_signal_214, sbe_n12}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U38 ( .a ({X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_217, sbe_Y_4_}), .c ({new_AGEMA_signal_222, sbe_n24}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U37 ( .a ({new_AGEMA_signal_203, sbe_Y_2_}), .b ({new_AGEMA_signal_209, sbe_n10}), .c ({new_AGEMA_signal_215, sbe_n23}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U36 ( .a ({new_AGEMA_signal_204, sbe_n9}), .b ({new_AGEMA_signal_197, sbe_n8}), .c ({new_AGEMA_signal_207, sbe_n22}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U35 ( .a ({X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_198, sbe_n11}), .c ({new_AGEMA_signal_201, sbe_n21}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U29 ( .a ({X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_209, sbe_n10}), .c ({new_AGEMA_signal_216, sbe_Y_6_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U28 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_194, sbe_Y_5_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U27 ( .a ({X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_209, sbe_n10}), .c ({new_AGEMA_signal_217, sbe_Y_4_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U26 ( .a ({X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_204, sbe_n9}), .c ({new_AGEMA_signal_209, sbe_n10}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U25 ( .a ({X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_197, sbe_n8}), .c ({new_AGEMA_signal_203, sbe_Y_2_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U24 ( .a ({X_s1[5], X_s0[5]}), .b ({X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_197, sbe_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U23 ( .a ({X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_206, sbe_n7}), .c ({new_AGEMA_signal_210, sbe_Y_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U22 ( .a ({X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_218, sbe_B_6_}), .c ({new_AGEMA_signal_223, sbe_Y_0_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U8 ( .a ({X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_211, sbe_n25}), .c ({new_AGEMA_signal_218, sbe_B_6_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U7 ( .a ({X_s1[5], X_s0[5]}), .b ({new_AGEMA_signal_204, sbe_n9}), .c ({new_AGEMA_signal_211, sbe_n25}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U6 ( .a ({X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_200, sbe_n2}), .c ({new_AGEMA_signal_204, sbe_n9}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U5 ( .a ({new_AGEMA_signal_212, sbe_n3}), .b ({new_AGEMA_signal_198, sbe_n11}), .c ({new_AGEMA_signal_219, sbe_B_3_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U4 ( .a ({X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_206, sbe_n7}), .c ({new_AGEMA_signal_212, sbe_n3}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U3 ( .a ({X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_200, sbe_n2}), .c ({new_AGEMA_signal_206, sbe_n7}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U2 ( .a ({X_s1[4], X_s0[4]}), .b ({X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_198, sbe_n11}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_U1 ( .a ({X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_200, sbe_n2}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m7_U2 ( .a ({new_AGEMA_signal_224, sbe_sel_in_m7_n8}), .b ({new_AGEMA_signal_230, sbe_Z[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_198, sbe_n11}), .a ({new_AGEMA_signal_215, sbe_n23}), .c ({new_AGEMA_signal_224, sbe_sel_in_m7_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m6_U2 ( .a ({new_AGEMA_signal_225, sbe_sel_in_m6_n8}), .b ({new_AGEMA_signal_231, sbe_Z[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_216, sbe_Y_6_}), .a ({new_AGEMA_signal_218, sbe_B_6_}), .c ({new_AGEMA_signal_225, sbe_sel_in_m6_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m5_U2 ( .a ({new_AGEMA_signal_226, sbe_sel_in_m5_n8}), .b ({new_AGEMA_signal_232, sbe_Z[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_194, sbe_Y_5_}), .a ({new_AGEMA_signal_214, sbe_n12}), .c ({new_AGEMA_signal_226, sbe_sel_in_m5_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m4_U2 ( .a ({new_AGEMA_signal_227, sbe_sel_in_m4_n8}), .b ({new_AGEMA_signal_233, sbe_Z[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_217, sbe_Y_4_}), .a ({new_AGEMA_signal_207, sbe_n22}), .c ({new_AGEMA_signal_227, sbe_sel_in_m4_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m3_U2 ( .a ({new_AGEMA_signal_228, sbe_sel_in_m3_n8}), .b ({new_AGEMA_signal_234, sbe_Z[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_201, sbe_n21}), .a ({new_AGEMA_signal_219, sbe_B_3_}), .c ({new_AGEMA_signal_228, sbe_sel_in_m3_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m2_U2 ( .a ({new_AGEMA_signal_213, sbe_sel_in_m2_n8}), .b ({new_AGEMA_signal_220, sbe_Z[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_203, sbe_Y_2_}), .a ({new_AGEMA_signal_200, sbe_n2}), .c ({new_AGEMA_signal_213, sbe_sel_in_m2_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m1_U2 ( .a ({new_AGEMA_signal_221, sbe_sel_in_m1_n8}), .b ({new_AGEMA_signal_229, sbe_Z[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_210, sbe_Y_1_}), .a ({new_AGEMA_signal_211, sbe_n25}), .c ({new_AGEMA_signal_221, sbe_sel_in_m1_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m0_U2 ( .a ({new_AGEMA_signal_235, sbe_sel_in_m0_n8}), .b ({new_AGEMA_signal_236, sbe_Z[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_in_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_223, sbe_Y_0_}), .a ({new_AGEMA_signal_222, sbe_n24}), .c ({new_AGEMA_signal_235, sbe_sel_in_m0_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U10 ( .a ({new_AGEMA_signal_236, sbe_Z[0]}), .b ({new_AGEMA_signal_229, sbe_Z[1]}), .c ({new_AGEMA_signal_250, sbe_inv_bl}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U9 ( .a ({new_AGEMA_signal_220, sbe_Z[2]}), .b ({new_AGEMA_signal_234, sbe_Z[3]}), .c ({new_AGEMA_signal_240, sbe_inv_bh}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U8 ( .a ({new_AGEMA_signal_251, sbe_inv_sb_0_}), .b ({new_AGEMA_signal_241, sbe_inv_sb_1_}), .c ({new_AGEMA_signal_258, sbe_inv_bb}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U7 ( .a ({new_AGEMA_signal_236, sbe_Z[0]}), .b ({new_AGEMA_signal_220, sbe_Z[2]}), .c ({new_AGEMA_signal_251, sbe_inv_sb_0_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U6 ( .a ({new_AGEMA_signal_234, sbe_Z[3]}), .b ({new_AGEMA_signal_229, sbe_Z[1]}), .c ({new_AGEMA_signal_241, sbe_inv_sb_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U5 ( .a ({new_AGEMA_signal_233, sbe_Z[4]}), .b ({new_AGEMA_signal_232, sbe_Z[5]}), .c ({new_AGEMA_signal_242, sbe_inv_al}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U4 ( .a ({new_AGEMA_signal_231, sbe_Z[6]}), .b ({new_AGEMA_signal_230, sbe_Z[7]}), .c ({new_AGEMA_signal_243, sbe_inv_ah}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U3 ( .a ({new_AGEMA_signal_244, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_245, sbe_inv_sa_1_}), .c ({new_AGEMA_signal_252, sbe_inv_aa}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U2 ( .a ({new_AGEMA_signal_233, sbe_Z[4]}), .b ({new_AGEMA_signal_231, sbe_Z[6]}), .c ({new_AGEMA_signal_244, sbe_inv_sa_0_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U1 ( .a ({new_AGEMA_signal_230, sbe_Z[7]}), .b ({new_AGEMA_signal_232, sbe_Z[5]}), .c ({new_AGEMA_signal_245, sbe_inv_sa_1_}) ) ;

    /* cells in depth 1 */
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U34 ( .a ({new_AGEMA_signal_264, sbe_inv_n21}), .b ({new_AGEMA_signal_259, sbe_inv_n20}), .c ({new_AGEMA_signal_268, sbe_inv_c[3]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U33 ( .a ({new_AGEMA_signal_253, sbe_inv_n19}), .b ({new_AGEMA_signal_237, sbe_inv_n18}), .c ({new_AGEMA_signal_259, sbe_inv_n20}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U32 ( .a ({new_AGEMA_signal_230, sbe_Z[7]}), .b ({new_AGEMA_signal_234, sbe_Z[3]}), .clk ( clk ), .r ({Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_237, sbe_inv_n18}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U31 ( .a ({new_AGEMA_signal_244, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_251, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[7], Fresh[6], Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_253, sbe_inv_n19}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U30 ( .a ({new_AGEMA_signal_262, sbe_inv_n17}), .b ({new_AGEMA_signal_247, sbe_inv_n16}), .c ({new_AGEMA_signal_264, sbe_inv_n21}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U29 ( .a ({new_AGEMA_signal_260, sbe_inv_n15}), .b ({new_AGEMA_signal_254, sbe_inv_n14}), .c ({new_AGEMA_signal_265, sbe_inv_c[2]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U28 ( .a ({new_AGEMA_signal_246, sbe_inv_n13}), .b ({new_AGEMA_signal_238, sbe_inv_n12}), .c ({new_AGEMA_signal_254, sbe_inv_n14}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U27 ( .a ({new_AGEMA_signal_231, sbe_Z[6]}), .b ({new_AGEMA_signal_220, sbe_Z[2]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_238, sbe_inv_n12}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U26 ( .a ({new_AGEMA_signal_245, sbe_inv_sa_1_}), .b ({new_AGEMA_signal_241, sbe_inv_sb_1_}), .clk ( clk ), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_246, sbe_inv_n13}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U25 ( .a ({new_AGEMA_signal_257, sbe_inv_n11}), .b ({new_AGEMA_signal_247, sbe_inv_n16}), .c ({new_AGEMA_signal_260, sbe_inv_n15}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U24 ( .a ({new_AGEMA_signal_243, sbe_inv_ah}), .b ({new_AGEMA_signal_240, sbe_inv_bh}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_247, sbe_inv_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U23 ( .a ({new_AGEMA_signal_266, sbe_inv_n10}), .b ({new_AGEMA_signal_261, sbe_inv_n9}), .c ({new_AGEMA_signal_269, sbe_inv_c[1]}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U22 ( .a ({new_AGEMA_signal_255, sbe_inv_n8}), .b ({new_AGEMA_signal_239, sbe_inv_n7}), .c ({new_AGEMA_signal_261, sbe_inv_n9}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U21 ( .a ({new_AGEMA_signal_229, sbe_Z[1]}), .b ({new_AGEMA_signal_232, sbe_Z[5]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_239, sbe_inv_n7}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U20 ( .a ({new_AGEMA_signal_242, sbe_inv_al}), .b ({new_AGEMA_signal_250, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_255, sbe_inv_n8}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U19 ( .a ({new_AGEMA_signal_262, sbe_inv_n17}), .b ({new_AGEMA_signal_257, sbe_inv_n11}), .c ({new_AGEMA_signal_266, sbe_inv_n10}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U18 ( .a ({new_AGEMA_signal_252, sbe_inv_aa}), .b ({new_AGEMA_signal_258, sbe_inv_bb}), .clk ( clk ), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_262, sbe_inv_n17}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U17 ( .a ({new_AGEMA_signal_257, sbe_inv_n11}), .b ({new_AGEMA_signal_267, sbe_inv_n6}), .c ({new_AGEMA_signal_270, sbe_inv_c[0]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U16 ( .a ({new_AGEMA_signal_249, sbe_inv_n5}), .b ({new_AGEMA_signal_263, sbe_inv_n4}), .c ({new_AGEMA_signal_267, sbe_inv_n6}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U15 ( .a ({new_AGEMA_signal_248, sbe_inv_n3}), .b ({new_AGEMA_signal_256, sbe_inv_n2}), .c ({new_AGEMA_signal_263, sbe_inv_n4}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U14 ( .a ({new_AGEMA_signal_242, sbe_inv_al}), .b ({new_AGEMA_signal_250, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_256, sbe_inv_n2}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U13 ( .a ({new_AGEMA_signal_233, sbe_Z[4]}), .b ({new_AGEMA_signal_236, sbe_Z[0]}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_248, sbe_inv_n3}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U12 ( .a ({new_AGEMA_signal_241, sbe_inv_sb_1_}), .b ({new_AGEMA_signal_245, sbe_inv_sa_1_}), .clk ( clk ), .r ({Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_249, sbe_inv_n5}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U11 ( .a ({new_AGEMA_signal_244, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_251, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_257, sbe_inv_n11}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U2 ( .a ({new_AGEMA_signal_265, sbe_inv_c[2]}), .b ({new_AGEMA_signal_268, sbe_inv_c[3]}), .c ({new_AGEMA_signal_273, sbe_inv_dinv_sa}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U1 ( .a ({new_AGEMA_signal_270, sbe_inv_c[0]}), .b ({new_AGEMA_signal_269, sbe_inv_c[1]}), .c ({new_AGEMA_signal_274, sbe_inv_dinv_sb}) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( sbe_Z[3] ), .Q ( new_AGEMA_signal_548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C ( clk ), .D ( new_AGEMA_signal_234 ), .Q ( new_AGEMA_signal_551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C ( clk ), .D ( sbe_Z[2] ), .Q ( new_AGEMA_signal_554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C ( clk ), .D ( new_AGEMA_signal_220 ), .Q ( new_AGEMA_signal_557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C ( clk ), .D ( sbe_inv_bh ), .Q ( new_AGEMA_signal_560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C ( clk ), .D ( new_AGEMA_signal_240 ), .Q ( new_AGEMA_signal_563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C ( clk ), .D ( sbe_Z[1] ), .Q ( new_AGEMA_signal_566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C ( clk ), .D ( new_AGEMA_signal_229 ), .Q ( new_AGEMA_signal_569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C ( clk ), .D ( sbe_Z[0] ), .Q ( new_AGEMA_signal_572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C ( clk ), .D ( new_AGEMA_signal_236 ), .Q ( new_AGEMA_signal_575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C ( clk ), .D ( sbe_inv_bl ), .Q ( new_AGEMA_signal_578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C ( clk ), .D ( new_AGEMA_signal_250 ), .Q ( new_AGEMA_signal_581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C ( clk ), .D ( sbe_inv_bb ), .Q ( new_AGEMA_signal_584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C ( clk ), .D ( new_AGEMA_signal_258 ), .Q ( new_AGEMA_signal_587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C ( clk ), .D ( sbe_inv_sb_1_ ), .Q ( new_AGEMA_signal_590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C ( clk ), .D ( new_AGEMA_signal_241 ), .Q ( new_AGEMA_signal_593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C ( clk ), .D ( sbe_inv_sb_0_ ), .Q ( new_AGEMA_signal_596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C ( clk ), .D ( new_AGEMA_signal_251 ), .Q ( new_AGEMA_signal_599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C ( clk ), .D ( sbe_Z[7] ), .Q ( new_AGEMA_signal_602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C ( clk ), .D ( new_AGEMA_signal_230 ), .Q ( new_AGEMA_signal_605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C ( clk ), .D ( sbe_Z[6] ), .Q ( new_AGEMA_signal_608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C ( clk ), .D ( new_AGEMA_signal_231 ), .Q ( new_AGEMA_signal_611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C ( clk ), .D ( sbe_inv_ah ), .Q ( new_AGEMA_signal_614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C ( clk ), .D ( new_AGEMA_signal_243 ), .Q ( new_AGEMA_signal_617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C ( clk ), .D ( sbe_Z[5] ), .Q ( new_AGEMA_signal_620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C ( clk ), .D ( new_AGEMA_signal_232 ), .Q ( new_AGEMA_signal_623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C ( clk ), .D ( sbe_Z[4] ), .Q ( new_AGEMA_signal_626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C ( clk ), .D ( new_AGEMA_signal_233 ), .Q ( new_AGEMA_signal_629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C ( clk ), .D ( sbe_inv_al ), .Q ( new_AGEMA_signal_632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C ( clk ), .D ( new_AGEMA_signal_242 ), .Q ( new_AGEMA_signal_635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C ( clk ), .D ( sbe_inv_aa ), .Q ( new_AGEMA_signal_638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C ( clk ), .D ( new_AGEMA_signal_252 ), .Q ( new_AGEMA_signal_641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C ( clk ), .D ( sbe_inv_sa_1_ ), .Q ( new_AGEMA_signal_644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C ( clk ), .D ( new_AGEMA_signal_245 ), .Q ( new_AGEMA_signal_647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C ( clk ), .D ( sbe_inv_sa_0_ ), .Q ( new_AGEMA_signal_650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C ( clk ), .D ( new_AGEMA_signal_244 ), .Q ( new_AGEMA_signal_653 ) ) ;

    /* cells in depth 2 */
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U9 ( .a ({new_AGEMA_signal_277, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_278, sbe_inv_dinv_d_1_}), .c ({new_AGEMA_signal_279, sbe_inv_dinv_sd}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U8 ( .a ({new_AGEMA_signal_271, sbe_inv_dinv_n4}), .b ({new_AGEMA_signal_275, sbe_inv_dinv_n3}), .c ({new_AGEMA_signal_277, sbe_inv_dinv_d_0_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U7 ( .a ({new_AGEMA_signal_274, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_273, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_275, sbe_inv_dinv_n3}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U6 ( .a ({new_AGEMA_signal_269, sbe_inv_c[1]}), .b ({new_AGEMA_signal_268, sbe_inv_c[3]}), .clk ( clk ), .r ({Fresh[55], Fresh[54], Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_271, sbe_inv_dinv_n4}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U5 ( .a ({new_AGEMA_signal_276, sbe_inv_dinv_n2}), .b ({new_AGEMA_signal_272, sbe_inv_dinv_n1}), .c ({new_AGEMA_signal_278, sbe_inv_dinv_d_1_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U4 ( .a ({new_AGEMA_signal_270, sbe_inv_c[0]}), .b ({new_AGEMA_signal_265, sbe_inv_c[2]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_272, sbe_inv_dinv_n1}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_U3 ( .a ({new_AGEMA_signal_274, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_273, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_276, sbe_inv_dinv_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( sbe_inv_c[1] ), .Q ( new_AGEMA_signal_536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_269 ), .Q ( new_AGEMA_signal_537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( sbe_inv_c[0] ), .Q ( new_AGEMA_signal_538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_270 ), .Q ( new_AGEMA_signal_539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( sbe_inv_dinv_sb ), .Q ( new_AGEMA_signal_540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_274 ), .Q ( new_AGEMA_signal_541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( sbe_inv_c[3] ), .Q ( new_AGEMA_signal_542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_268 ), .Q ( new_AGEMA_signal_543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( sbe_inv_c[2] ), .Q ( new_AGEMA_signal_544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_265 ), .Q ( new_AGEMA_signal_545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( sbe_inv_dinv_sa ), .Q ( new_AGEMA_signal_546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_273 ), .Q ( new_AGEMA_signal_547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_548 ), .Q ( new_AGEMA_signal_549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C ( clk ), .D ( new_AGEMA_signal_551 ), .Q ( new_AGEMA_signal_552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C ( clk ), .D ( new_AGEMA_signal_554 ), .Q ( new_AGEMA_signal_555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C ( clk ), .D ( new_AGEMA_signal_557 ), .Q ( new_AGEMA_signal_558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C ( clk ), .D ( new_AGEMA_signal_560 ), .Q ( new_AGEMA_signal_561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C ( clk ), .D ( new_AGEMA_signal_563 ), .Q ( new_AGEMA_signal_564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C ( clk ), .D ( new_AGEMA_signal_566 ), .Q ( new_AGEMA_signal_567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C ( clk ), .D ( new_AGEMA_signal_569 ), .Q ( new_AGEMA_signal_570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C ( clk ), .D ( new_AGEMA_signal_572 ), .Q ( new_AGEMA_signal_573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C ( clk ), .D ( new_AGEMA_signal_575 ), .Q ( new_AGEMA_signal_576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C ( clk ), .D ( new_AGEMA_signal_578 ), .Q ( new_AGEMA_signal_579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C ( clk ), .D ( new_AGEMA_signal_581 ), .Q ( new_AGEMA_signal_582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C ( clk ), .D ( new_AGEMA_signal_584 ), .Q ( new_AGEMA_signal_585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C ( clk ), .D ( new_AGEMA_signal_587 ), .Q ( new_AGEMA_signal_588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C ( clk ), .D ( new_AGEMA_signal_590 ), .Q ( new_AGEMA_signal_591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C ( clk ), .D ( new_AGEMA_signal_593 ), .Q ( new_AGEMA_signal_594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C ( clk ), .D ( new_AGEMA_signal_596 ), .Q ( new_AGEMA_signal_597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C ( clk ), .D ( new_AGEMA_signal_599 ), .Q ( new_AGEMA_signal_600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C ( clk ), .D ( new_AGEMA_signal_602 ), .Q ( new_AGEMA_signal_603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C ( clk ), .D ( new_AGEMA_signal_605 ), .Q ( new_AGEMA_signal_606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C ( clk ), .D ( new_AGEMA_signal_608 ), .Q ( new_AGEMA_signal_609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C ( clk ), .D ( new_AGEMA_signal_611 ), .Q ( new_AGEMA_signal_612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C ( clk ), .D ( new_AGEMA_signal_614 ), .Q ( new_AGEMA_signal_615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C ( clk ), .D ( new_AGEMA_signal_617 ), .Q ( new_AGEMA_signal_618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C ( clk ), .D ( new_AGEMA_signal_620 ), .Q ( new_AGEMA_signal_621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C ( clk ), .D ( new_AGEMA_signal_623 ), .Q ( new_AGEMA_signal_624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C ( clk ), .D ( new_AGEMA_signal_626 ), .Q ( new_AGEMA_signal_627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C ( clk ), .D ( new_AGEMA_signal_629 ), .Q ( new_AGEMA_signal_630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C ( clk ), .D ( new_AGEMA_signal_632 ), .Q ( new_AGEMA_signal_633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C ( clk ), .D ( new_AGEMA_signal_635 ), .Q ( new_AGEMA_signal_636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C ( clk ), .D ( new_AGEMA_signal_638 ), .Q ( new_AGEMA_signal_639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C ( clk ), .D ( new_AGEMA_signal_641 ), .Q ( new_AGEMA_signal_642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C ( clk ), .D ( new_AGEMA_signal_644 ), .Q ( new_AGEMA_signal_645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C ( clk ), .D ( new_AGEMA_signal_647 ), .Q ( new_AGEMA_signal_648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C ( clk ), .D ( new_AGEMA_signal_650 ), .Q ( new_AGEMA_signal_651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C ( clk ), .D ( new_AGEMA_signal_653 ), .Q ( new_AGEMA_signal_654 ) ) ;

    /* cells in depth 3 */
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U39 ( .a ({new_AGEMA_signal_289, sbe_inv_d_0_}), .b ({new_AGEMA_signal_288, sbe_inv_d_1_}), .c ({new_AGEMA_signal_290, sbe_inv_dl}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U38 ( .a ({new_AGEMA_signal_287, sbe_inv_d_2_}), .b ({new_AGEMA_signal_286, sbe_inv_d_3_}), .c ({new_AGEMA_signal_291, sbe_inv_dh}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U37 ( .a ({new_AGEMA_signal_292, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_293, sbe_inv_sd_1_}), .c ({new_AGEMA_signal_302, sbe_inv_dd}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U36 ( .a ({new_AGEMA_signal_289, sbe_inv_d_0_}), .b ({new_AGEMA_signal_287, sbe_inv_d_2_}), .c ({new_AGEMA_signal_292, sbe_inv_sd_0_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_U35 ( .a ({new_AGEMA_signal_288, sbe_inv_d_1_}), .b ({new_AGEMA_signal_286, sbe_inv_d_3_}), .c ({new_AGEMA_signal_293, sbe_inv_sd_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_pmul_U5 ( .a ({new_AGEMA_signal_284, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_280, sbe_inv_dinv_pmul_n8}), .c ({new_AGEMA_signal_286, sbe_inv_d_3_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_pmul_U4 ( .a ({new_AGEMA_signal_278, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_537, new_AGEMA_signal_536}), .clk ( clk ), .r ({Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_280, sbe_inv_dinv_pmul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_pmul_U3 ( .a ({new_AGEMA_signal_284, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_281, sbe_inv_dinv_pmul_n7}), .c ({new_AGEMA_signal_287, sbe_inv_d_2_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_pmul_U2 ( .a ({new_AGEMA_signal_277, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_539, new_AGEMA_signal_538}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_281, sbe_inv_dinv_pmul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_pmul_U1 ( .a ({new_AGEMA_signal_279, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_541, new_AGEMA_signal_540}), .clk ( clk ), .r ({Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_284, sbe_inv_dinv_pmul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_qmul_U5 ( .a ({new_AGEMA_signal_285, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_282, sbe_inv_dinv_qmul_n8}), .c ({new_AGEMA_signal_288, sbe_inv_d_1_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_qmul_U4 ( .a ({new_AGEMA_signal_278, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_543, new_AGEMA_signal_542}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_282, sbe_inv_dinv_qmul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_qmul_U3 ( .a ({new_AGEMA_signal_285, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_283, sbe_inv_dinv_qmul_n7}), .c ({new_AGEMA_signal_289, sbe_inv_d_0_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_qmul_U2 ( .a ({new_AGEMA_signal_277, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_545, new_AGEMA_signal_544}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_283, sbe_inv_dinv_qmul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_dinv_qmul_U1 ( .a ({new_AGEMA_signal_279, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_547, new_AGEMA_signal_546}), .clk ( clk ), .r ({Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_285, sbe_inv_dinv_qmul_n9}) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_549 ), .Q ( new_AGEMA_signal_550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C ( clk ), .D ( new_AGEMA_signal_552 ), .Q ( new_AGEMA_signal_553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C ( clk ), .D ( new_AGEMA_signal_555 ), .Q ( new_AGEMA_signal_556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C ( clk ), .D ( new_AGEMA_signal_558 ), .Q ( new_AGEMA_signal_559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C ( clk ), .D ( new_AGEMA_signal_561 ), .Q ( new_AGEMA_signal_562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C ( clk ), .D ( new_AGEMA_signal_564 ), .Q ( new_AGEMA_signal_565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C ( clk ), .D ( new_AGEMA_signal_567 ), .Q ( new_AGEMA_signal_568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C ( clk ), .D ( new_AGEMA_signal_570 ), .Q ( new_AGEMA_signal_571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C ( clk ), .D ( new_AGEMA_signal_573 ), .Q ( new_AGEMA_signal_574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C ( clk ), .D ( new_AGEMA_signal_576 ), .Q ( new_AGEMA_signal_577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C ( clk ), .D ( new_AGEMA_signal_579 ), .Q ( new_AGEMA_signal_580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C ( clk ), .D ( new_AGEMA_signal_582 ), .Q ( new_AGEMA_signal_583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C ( clk ), .D ( new_AGEMA_signal_585 ), .Q ( new_AGEMA_signal_586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C ( clk ), .D ( new_AGEMA_signal_588 ), .Q ( new_AGEMA_signal_589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C ( clk ), .D ( new_AGEMA_signal_591 ), .Q ( new_AGEMA_signal_592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C ( clk ), .D ( new_AGEMA_signal_594 ), .Q ( new_AGEMA_signal_595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C ( clk ), .D ( new_AGEMA_signal_597 ), .Q ( new_AGEMA_signal_598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C ( clk ), .D ( new_AGEMA_signal_600 ), .Q ( new_AGEMA_signal_601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C ( clk ), .D ( new_AGEMA_signal_603 ), .Q ( new_AGEMA_signal_604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C ( clk ), .D ( new_AGEMA_signal_606 ), .Q ( new_AGEMA_signal_607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C ( clk ), .D ( new_AGEMA_signal_609 ), .Q ( new_AGEMA_signal_610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C ( clk ), .D ( new_AGEMA_signal_612 ), .Q ( new_AGEMA_signal_613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C ( clk ), .D ( new_AGEMA_signal_615 ), .Q ( new_AGEMA_signal_616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C ( clk ), .D ( new_AGEMA_signal_618 ), .Q ( new_AGEMA_signal_619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C ( clk ), .D ( new_AGEMA_signal_621 ), .Q ( new_AGEMA_signal_622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C ( clk ), .D ( new_AGEMA_signal_624 ), .Q ( new_AGEMA_signal_625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C ( clk ), .D ( new_AGEMA_signal_627 ), .Q ( new_AGEMA_signal_628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C ( clk ), .D ( new_AGEMA_signal_630 ), .Q ( new_AGEMA_signal_631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C ( clk ), .D ( new_AGEMA_signal_633 ), .Q ( new_AGEMA_signal_634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C ( clk ), .D ( new_AGEMA_signal_636 ), .Q ( new_AGEMA_signal_637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C ( clk ), .D ( new_AGEMA_signal_639 ), .Q ( new_AGEMA_signal_640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C ( clk ), .D ( new_AGEMA_signal_642 ), .Q ( new_AGEMA_signal_643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C ( clk ), .D ( new_AGEMA_signal_645 ), .Q ( new_AGEMA_signal_646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C ( clk ), .D ( new_AGEMA_signal_648 ), .Q ( new_AGEMA_signal_649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C ( clk ), .D ( new_AGEMA_signal_651 ), .Q ( new_AGEMA_signal_652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C ( clk ), .D ( new_AGEMA_signal_654 ), .Q ( new_AGEMA_signal_655 ) ) ;

    /* cells in depth 4 */
    not_masked #(.low_latency(1), .pipeline(1)) sbe_U40 ( .a ({new_AGEMA_signal_326, sbe_C_2_}), .b ({new_AGEMA_signal_329, sbe_n1}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U34 ( .a ({new_AGEMA_signal_332, sbe_C_7_}), .b ({new_AGEMA_signal_342, sbe_n17}), .c ({new_AGEMA_signal_347, sbe_n16}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U33 ( .a ({new_AGEMA_signal_324, sbe_C_4_}), .b ({new_AGEMA_signal_336, sbe_n18}), .c ({new_AGEMA_signal_342, sbe_n17}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U32 ( .a ({new_AGEMA_signal_333, sbe_C_5_}), .b ({new_AGEMA_signal_335, sbe_C_1_}), .c ({new_AGEMA_signal_336, sbe_n18}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U31 ( .a ({new_AGEMA_signal_335, sbe_C_1_}), .b ({new_AGEMA_signal_324, sbe_C_4_}), .c ({new_AGEMA_signal_337, sbe_n15}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U30 ( .a ({new_AGEMA_signal_323, sbe_C_6_}), .b ({new_AGEMA_signal_335, sbe_C_1_}), .c ({new_AGEMA_signal_338, sbe_n14}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U21 ( .a ({new_AGEMA_signal_348, sbe_n6}), .b ({new_AGEMA_signal_335, sbe_C_1_}), .c ({new_AGEMA_signal_356, sbe_X[6]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U20 ( .a ({new_AGEMA_signal_326, sbe_C_2_}), .b ({new_AGEMA_signal_348, sbe_n6}), .c ({new_AGEMA_signal_357, sbe_X[5]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U19 ( .a ({new_AGEMA_signal_330, sbe_D_5_}), .b ({new_AGEMA_signal_343, sbe_n20}), .c ({new_AGEMA_signal_348, sbe_n6}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U18 ( .a ({new_AGEMA_signal_344, sbe_n5}), .b ({new_AGEMA_signal_341, sbe_D_0_}), .c ({new_AGEMA_signal_349, sbe_X[3]}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U17 ( .a ({new_AGEMA_signal_343, sbe_n20}), .b ({new_AGEMA_signal_331, sbe_n4}), .c ({new_AGEMA_signal_350, sbe_D_3_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U16 ( .a ({new_AGEMA_signal_333, sbe_C_5_}), .b ({new_AGEMA_signal_339, sbe_D_6_}), .c ({new_AGEMA_signal_343, sbe_n20}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U15 ( .a ({new_AGEMA_signal_332, sbe_C_7_}), .b ({new_AGEMA_signal_334, sbe_C_3_}), .c ({new_AGEMA_signal_339, sbe_D_6_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U14 ( .a ({new_AGEMA_signal_330, sbe_D_5_}), .b ({new_AGEMA_signal_344, sbe_n5}), .c ({new_AGEMA_signal_351, sbe_D_2_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U13 ( .a ({new_AGEMA_signal_326, sbe_C_2_}), .b ({new_AGEMA_signal_340, sbe_n19}), .c ({new_AGEMA_signal_344, sbe_n5}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U12 ( .a ({new_AGEMA_signal_333, sbe_C_5_}), .b ({new_AGEMA_signal_334, sbe_C_3_}), .c ({new_AGEMA_signal_340, sbe_n19}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U11 ( .a ({new_AGEMA_signal_323, sbe_C_6_}), .b ({new_AGEMA_signal_327, sbe_C_0_}), .c ({new_AGEMA_signal_330, sbe_D_5_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U10 ( .a ({new_AGEMA_signal_335, sbe_C_1_}), .b ({new_AGEMA_signal_331, sbe_n4}), .c ({new_AGEMA_signal_341, sbe_D_0_}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) sbe_U9 ( .a ({new_AGEMA_signal_323, sbe_C_6_}), .b ({new_AGEMA_signal_324, sbe_C_4_}), .c ({new_AGEMA_signal_331, sbe_n4}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_U4 ( .a ({new_AGEMA_signal_325, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_311, sbe_inv_pmul_ph[1]}), .c ({new_AGEMA_signal_332, sbe_C_7_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_U3 ( .a ({new_AGEMA_signal_316, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_312, sbe_inv_pmul_ph[0]}), .c ({new_AGEMA_signal_323, sbe_C_6_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_U2 ( .a ({new_AGEMA_signal_325, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_313, sbe_inv_pmul_pl[1]}), .c ({new_AGEMA_signal_333, sbe_C_5_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_U1 ( .a ({new_AGEMA_signal_316, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_314, sbe_inv_pmul_pl[0]}), .c ({new_AGEMA_signal_324, sbe_C_4_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_himul_U5 ( .a ({new_AGEMA_signal_303, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_294, sbe_inv_pmul_himul_n8}), .c ({new_AGEMA_signal_311, sbe_inv_pmul_ph[1]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_himul_U4 ( .a ({new_AGEMA_signal_286, sbe_inv_d_3_}), .b ({new_AGEMA_signal_553, new_AGEMA_signal_550}), .clk ( clk ), .r ({Fresh[91], Fresh[90], Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_294, sbe_inv_pmul_himul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_himul_U3 ( .a ({new_AGEMA_signal_303, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_295, sbe_inv_pmul_himul_n7}), .c ({new_AGEMA_signal_312, sbe_inv_pmul_ph[0]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_himul_U2 ( .a ({new_AGEMA_signal_287, sbe_inv_d_2_}), .b ({new_AGEMA_signal_559, new_AGEMA_signal_556}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_295, sbe_inv_pmul_himul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_himul_U1 ( .a ({new_AGEMA_signal_291, sbe_inv_dh}), .b ({new_AGEMA_signal_565, new_AGEMA_signal_562}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_303, sbe_inv_pmul_himul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_lomul_U5 ( .a ({new_AGEMA_signal_304, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_296, sbe_inv_pmul_lomul_n8}), .c ({new_AGEMA_signal_313, sbe_inv_pmul_pl[1]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_lomul_U4 ( .a ({new_AGEMA_signal_288, sbe_inv_d_1_}), .b ({new_AGEMA_signal_571, new_AGEMA_signal_568}), .clk ( clk ), .r ({Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_296, sbe_inv_pmul_lomul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_lomul_U3 ( .a ({new_AGEMA_signal_304, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_297, sbe_inv_pmul_lomul_n7}), .c ({new_AGEMA_signal_314, sbe_inv_pmul_pl[0]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_lomul_U2 ( .a ({new_AGEMA_signal_289, sbe_inv_d_0_}), .b ({new_AGEMA_signal_577, new_AGEMA_signal_574}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_297, sbe_inv_pmul_lomul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_lomul_U1 ( .a ({new_AGEMA_signal_290, sbe_inv_dl}), .b ({new_AGEMA_signal_583, new_AGEMA_signal_580}), .clk ( clk ), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_304, sbe_inv_pmul_lomul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_summul_U5 ( .a ({new_AGEMA_signal_306, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_315, sbe_inv_pmul_summul_n8}), .c ({new_AGEMA_signal_325, sbe_inv_pmul_p_1_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_summul_U4 ( .a ({new_AGEMA_signal_302, sbe_inv_dd}), .b ({new_AGEMA_signal_589, new_AGEMA_signal_586}), .clk ( clk ), .r ({Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_315, sbe_inv_pmul_summul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_summul_U3 ( .a ({new_AGEMA_signal_306, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_305, sbe_inv_pmul_summul_n7}), .c ({new_AGEMA_signal_316, sbe_inv_pmul_p_0_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_summul_U2 ( .a ({new_AGEMA_signal_293, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_595, new_AGEMA_signal_592}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_305, sbe_inv_pmul_summul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_pmul_summul_U1 ( .a ({new_AGEMA_signal_292, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_601, new_AGEMA_signal_598}), .clk ( clk ), .r ({Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_306, sbe_inv_pmul_summul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_U4 ( .a ({new_AGEMA_signal_328, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_317, sbe_inv_qmul_ph[1]}), .c ({new_AGEMA_signal_334, sbe_C_3_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_U3 ( .a ({new_AGEMA_signal_322, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_318, sbe_inv_qmul_ph[0]}), .c ({new_AGEMA_signal_326, sbe_C_2_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_U2 ( .a ({new_AGEMA_signal_328, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_319, sbe_inv_qmul_pl[1]}), .c ({new_AGEMA_signal_335, sbe_C_1_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_U1 ( .a ({new_AGEMA_signal_322, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_320, sbe_inv_qmul_pl[0]}), .c ({new_AGEMA_signal_327, sbe_C_0_}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_himul_U5 ( .a ({new_AGEMA_signal_307, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_298, sbe_inv_qmul_himul_n8}), .c ({new_AGEMA_signal_317, sbe_inv_qmul_ph[1]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_himul_U4 ( .a ({new_AGEMA_signal_286, sbe_inv_d_3_}), .b ({new_AGEMA_signal_607, new_AGEMA_signal_604}), .clk ( clk ), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_298, sbe_inv_qmul_himul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_himul_U3 ( .a ({new_AGEMA_signal_307, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_299, sbe_inv_qmul_himul_n7}), .c ({new_AGEMA_signal_318, sbe_inv_qmul_ph[0]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_himul_U2 ( .a ({new_AGEMA_signal_287, sbe_inv_d_2_}), .b ({new_AGEMA_signal_613, new_AGEMA_signal_610}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_299, sbe_inv_qmul_himul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_himul_U1 ( .a ({new_AGEMA_signal_291, sbe_inv_dh}), .b ({new_AGEMA_signal_619, new_AGEMA_signal_616}), .clk ( clk ), .r ({Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_307, sbe_inv_qmul_himul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_lomul_U5 ( .a ({new_AGEMA_signal_308, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_300, sbe_inv_qmul_lomul_n8}), .c ({new_AGEMA_signal_319, sbe_inv_qmul_pl[1]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_lomul_U4 ( .a ({new_AGEMA_signal_288, sbe_inv_d_1_}), .b ({new_AGEMA_signal_625, new_AGEMA_signal_622}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136]}), .c ({new_AGEMA_signal_300, sbe_inv_qmul_lomul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_lomul_U3 ( .a ({new_AGEMA_signal_308, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_301, sbe_inv_qmul_lomul_n7}), .c ({new_AGEMA_signal_320, sbe_inv_qmul_pl[0]}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_lomul_U2 ( .a ({new_AGEMA_signal_289, sbe_inv_d_0_}), .b ({new_AGEMA_signal_631, new_AGEMA_signal_628}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_301, sbe_inv_qmul_lomul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_lomul_U1 ( .a ({new_AGEMA_signal_290, sbe_inv_dl}), .b ({new_AGEMA_signal_637, new_AGEMA_signal_634}), .clk ( clk ), .r ({Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_308, sbe_inv_qmul_lomul_n9}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_summul_U5 ( .a ({new_AGEMA_signal_310, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_321, sbe_inv_qmul_summul_n8}), .c ({new_AGEMA_signal_328, sbe_inv_qmul_p_1_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_summul_U4 ( .a ({new_AGEMA_signal_302, sbe_inv_dd}), .b ({new_AGEMA_signal_643, new_AGEMA_signal_640}), .clk ( clk ), .r ({Fresh[151], Fresh[150], Fresh[149], Fresh[148]}), .c ({new_AGEMA_signal_321, sbe_inv_qmul_summul_n8}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_summul_U3 ( .a ({new_AGEMA_signal_310, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_309, sbe_inv_qmul_summul_n7}), .c ({new_AGEMA_signal_322, sbe_inv_qmul_p_0_}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_summul_U2 ( .a ({new_AGEMA_signal_293, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_649, new_AGEMA_signal_646}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152]}), .c ({new_AGEMA_signal_309, sbe_inv_qmul_summul_n7}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) sbe_inv_qmul_summul_U1 ( .a ({new_AGEMA_signal_292, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_655, new_AGEMA_signal_652}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_310, sbe_inv_qmul_summul_n9}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m7_U2 ( .a ({new_AGEMA_signal_345, sbe_sel_out_m7_n8}), .b ({new_AGEMA_signal_352, O[7]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_337, sbe_n15}), .a ({new_AGEMA_signal_340, sbe_n19}), .c ({new_AGEMA_signal_345, sbe_sel_out_m7_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m6_U2 ( .a ({new_AGEMA_signal_362, sbe_sel_out_m6_n8}), .b ({new_AGEMA_signal_366, O[6]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_356, sbe_X[6]}), .a ({new_AGEMA_signal_339, sbe_D_6_}), .c ({new_AGEMA_signal_362, sbe_sel_out_m6_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m5_U2 ( .a ({new_AGEMA_signal_363, sbe_sel_out_m5_n8}), .b ({new_AGEMA_signal_367, O[5]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_357, sbe_X[5]}), .a ({new_AGEMA_signal_330, sbe_D_5_}), .c ({new_AGEMA_signal_363, sbe_sel_out_m5_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m4_U2 ( .a ({new_AGEMA_signal_353, sbe_sel_out_m4_n8}), .b ({new_AGEMA_signal_358, O[4]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_338, sbe_n14}), .a ({new_AGEMA_signal_343, sbe_n20}), .c ({new_AGEMA_signal_353, sbe_sel_out_m4_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m3_U2 ( .a ({new_AGEMA_signal_359, sbe_sel_out_m3_n8}), .b ({new_AGEMA_signal_364, O[3]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_349, sbe_X[3]}), .a ({new_AGEMA_signal_350, sbe_D_3_}), .c ({new_AGEMA_signal_359, sbe_sel_out_m3_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m2_U2 ( .a ({new_AGEMA_signal_360, sbe_sel_out_m2_n8}), .b ({new_AGEMA_signal_365, O[2]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_347, sbe_n16}), .a ({new_AGEMA_signal_351, sbe_D_2_}), .c ({new_AGEMA_signal_360, sbe_sel_out_m2_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m1_U2 ( .a ({new_AGEMA_signal_354, sbe_sel_out_m1_n8}), .b ({new_AGEMA_signal_361, O[1]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_336, sbe_n18}), .a ({new_AGEMA_signal_342, sbe_n17}), .c ({new_AGEMA_signal_354, sbe_sel_out_m1_n8}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m0_U2 ( .a ({new_AGEMA_signal_346, sbe_sel_out_m0_n8}), .b ({new_AGEMA_signal_355, O[0]}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) sbe_sel_out_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_329, sbe_n1}), .a ({new_AGEMA_signal_341, sbe_D_0_}), .c ({new_AGEMA_signal_346, sbe_sel_out_m0_n8}) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_352, O[7]}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_366, O[6]}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_367, O[5]}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_358, O[4]}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_364, O[3]}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_365, O[2]}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_361, O[1]}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) Y_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_355, O[0]}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
