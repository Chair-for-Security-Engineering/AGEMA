/* modified netlist. Source: module AES in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module AES_GHPC_ANF_ClockGating_d1 (plaintext_s0, key_s0, clk, start, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [7:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_677 ;
    wire signal_679 ;
    wire signal_681 ;
    wire signal_683 ;
    wire signal_685 ;
    wire signal_687 ;
    wire signal_689 ;
    wire signal_691 ;
    wire signal_693 ;
    wire signal_695 ;
    wire signal_697 ;
    wire signal_699 ;
    wire signal_701 ;
    wire signal_703 ;
    wire signal_705 ;
    wire signal_707 ;
    wire signal_709 ;
    wire signal_711 ;
    wire signal_713 ;
    wire signal_715 ;
    wire signal_717 ;
    wire signal_719 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2024 ;
    wire signal_2027 ;
    wire signal_2030 ;
    wire signal_2033 ;
    wire signal_2036 ;
    wire signal_2039 ;
    wire signal_2042 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2051 ;
    wire signal_2053 ;
    wire signal_2055 ;
    wire signal_2058 ;
    wire signal_2060 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2156 ;
    wire signal_2159 ;
    wire signal_2162 ;
    wire signal_2165 ;
    wire signal_2168 ;
    wire signal_2171 ;
    wire signal_2174 ;
    wire signal_2177 ;
    wire signal_2180 ;
    wire signal_2183 ;
    wire signal_2186 ;
    wire signal_2189 ;
    wire signal_2192 ;
    wire signal_2195 ;
    wire signal_2198 ;
    wire signal_2201 ;
    wire signal_2204 ;
    wire signal_2207 ;
    wire signal_2210 ;
    wire signal_2213 ;
    wire signal_2216 ;
    wire signal_2219 ;
    wire signal_2222 ;
    wire signal_2225 ;
    wire signal_2228 ;
    wire signal_2231 ;
    wire signal_2234 ;
    wire signal_2237 ;
    wire signal_2240 ;
    wire signal_2243 ;
    wire signal_2246 ;
    wire signal_2249 ;
    wire signal_2252 ;
    wire signal_2255 ;
    wire signal_2258 ;
    wire signal_2261 ;
    wire signal_2264 ;
    wire signal_2267 ;
    wire signal_2270 ;
    wire signal_2273 ;
    wire signal_2276 ;
    wire signal_2279 ;
    wire signal_2282 ;
    wire signal_2285 ;
    wire signal_2288 ;
    wire signal_2291 ;
    wire signal_2294 ;
    wire signal_2297 ;
    wire signal_2300 ;
    wire signal_2303 ;
    wire signal_2306 ;
    wire signal_2309 ;
    wire signal_2312 ;
    wire signal_2315 ;
    wire signal_2318 ;
    wire signal_2321 ;
    wire signal_2324 ;
    wire signal_2327 ;
    wire signal_2330 ;
    wire signal_2333 ;
    wire signal_2336 ;
    wire signal_2339 ;
    wire signal_2342 ;
    wire signal_2345 ;
    wire signal_2348 ;
    wire signal_2351 ;
    wire signal_2354 ;
    wire signal_2357 ;
    wire signal_2360 ;
    wire signal_2363 ;
    wire signal_2366 ;
    wire signal_2369 ;
    wire signal_2372 ;
    wire signal_2375 ;
    wire signal_2378 ;
    wire signal_2381 ;
    wire signal_2384 ;
    wire signal_2387 ;
    wire signal_2390 ;
    wire signal_2393 ;
    wire signal_2396 ;
    wire signal_2399 ;
    wire signal_2402 ;
    wire signal_2405 ;
    wire signal_2408 ;
    wire signal_2411 ;
    wire signal_2414 ;
    wire signal_2417 ;
    wire signal_2420 ;
    wire signal_2423 ;
    wire signal_2426 ;
    wire signal_2429 ;
    wire signal_2432 ;
    wire signal_2435 ;
    wire signal_2438 ;
    wire signal_2441 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2779 ;
    wire signal_2781 ;
    wire signal_2783 ;
    wire signal_2785 ;
    wire signal_2787 ;
    wire signal_2789 ;
    wire signal_2791 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3247 ;
    wire signal_3249 ;
    wire signal_3251 ;
    wire signal_3253 ;
    wire signal_3255 ;
    wire signal_3257 ;
    wire signal_3259 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3273 ;
    wire signal_3275 ;
    wire signal_3277 ;
    wire signal_3279 ;
    wire signal_3281 ;
    wire signal_3283 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3422 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_404) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_1983, signal_1493}), .c ({signal_1984, signal_1413}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_2 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_1986, signal_1492}), .c ({signal_1987, signal_1412}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_3 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_1989, signal_1491}), .c ({signal_1990, signal_1411}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_4 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_1992, signal_1490}), .c ({signal_1993, signal_1410}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_5 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_1995, signal_1489}), .c ({signal_1996, signal_1409}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_6 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_1998, signal_1488}), .c ({signal_1999, signal_1408}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_7 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2001, signal_1487}), .c ({signal_2002, signal_1407}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_8 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2004, signal_1486}), .c ({signal_2005, signal_1406}) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_399), .A2 (signal_398), .ZN (signal_405) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_402), .A2 (signal_405), .ZN (done) ) ;
    AND2_X1 cell_11 ( .A1 (signal_401), .A2 (signal_396), .ZN (signal_400) ) ;
    INV_X1 cell_12 ( .A (start), .ZN (signal_403) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_406), .A2 (signal_415), .ZN (signal_422) ) ;
    XNOR2_X1 cell_14 ( .A (signal_424), .B (signal_425), .ZN (signal_423) ) ;
    NOR2_X1 cell_15 ( .A1 (signal_407), .A2 (signal_408), .ZN (signal_398) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_421), .A2 (signal_416), .ZN (signal_408) ) ;
    INV_X1 cell_17 ( .A (signal_406), .ZN (signal_407) ) ;
    INV_X1 cell_18 ( .A (signal_420), .ZN (signal_416) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_409), .A2 (signal_410), .ZN (signal_419) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_396), .A2 (signal_418), .ZN (signal_409) ) ;
    NOR2_X1 cell_21 ( .A1 (signal_427), .A2 (signal_424), .ZN (signal_413) ) ;
    NOR2_X1 cell_22 ( .A1 (signal_425), .A2 (signal_428), .ZN (signal_412) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_415), .A2 (signal_414), .ZN (signal_396) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_414) ) ;
    INV_X1 cell_25 ( .A (signal_393), .ZN (signal_415) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_412), .A2 (signal_413), .ZN (signal_411) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_426), .A2 (signal_411), .ZN (signal_406) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_393), .A2 (signal_406), .ZN (signal_410) ) ;
    INV_X1 cell_29 ( .A (signal_410), .ZN (signal_395) ) ;
    NOR2_X1 cell_30 ( .A1 (signal_417), .A2 (signal_415), .ZN (signal_394) ) ;
    MUX2_X1 cell_31 ( .S (signal_393), .A (1'b1), .B (signal_423), .Z (signal_429) ) ;
    MUX2_X1 cell_34 ( .S (signal_393), .A (1'b0), .B (signal_425), .Z (signal_431) ) ;
    MUX2_X1 cell_37 ( .S (signal_393), .A (1'b1), .B (signal_426), .Z (signal_433) ) ;
    MUX2_X1 cell_40 ( .S (signal_393), .A (1'b0), .B (signal_427), .Z (signal_435) ) ;
    MUX2_X1 cell_43 ( .S (signal_393), .A (1'b1), .B (signal_428), .Z (signal_437) ) ;
    MUX2_X1 cell_46 ( .S (signal_422), .A (1'b1), .B (signal_416), .Z (signal_439) ) ;
    MUX2_X1 cell_49 ( .S (signal_422), .A (1'b0), .B (signal_421), .Z (signal_441) ) ;
    INV_X1 cell_52 ( .A (signal_418), .ZN (signal_417) ) ;
    INV_X1 cell_64 ( .A (signal_394), .ZN (signal_453) ) ;
    INV_X1 cell_65 ( .A (signal_453), .ZN (signal_455) ) ;
    INV_X1 cell_66 ( .A (signal_393), .ZN (signal_444) ) ;
    INV_X1 cell_67 ( .A (signal_444), .ZN (signal_452) ) ;
    INV_X1 cell_68 ( .A (signal_456), .ZN (signal_464) ) ;
    INV_X1 cell_69 ( .A (signal_453), .ZN (signal_454) ) ;
    INV_X1 cell_70 ( .A (signal_444), .ZN (signal_448) ) ;
    INV_X1 cell_71 ( .A (signal_456), .ZN (signal_460) ) ;
    INV_X1 cell_72 ( .A (signal_444), .ZN (signal_446) ) ;
    INV_X1 cell_73 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_74 ( .A (signal_444), .ZN (signal_450) ) ;
    INV_X1 cell_75 ( .A (signal_456), .ZN (signal_462) ) ;
    INV_X1 cell_76 ( .A (signal_444), .ZN (signal_445) ) ;
    INV_X1 cell_77 ( .A (signal_456), .ZN (signal_457) ) ;
    INV_X1 cell_78 ( .A (signal_444), .ZN (signal_447) ) ;
    INV_X1 cell_79 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_80 ( .A (signal_444), .ZN (signal_449) ) ;
    INV_X1 cell_81 ( .A (signal_456), .ZN (signal_461) ) ;
    INV_X1 cell_82 ( .A (signal_444), .ZN (signal_451) ) ;
    INV_X1 cell_83 ( .A (signal_456), .ZN (signal_463) ) ;
    INV_X1 cell_84 ( .A (signal_395), .ZN (signal_456) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_85 ( .s (signal_457), .b ({signal_2156, signal_1677}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_3126, signal_465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_88 ( .s (signal_457), .b ({signal_2159, signal_1676}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_3127, signal_467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_91 ( .s (signal_457), .b ({signal_2162, signal_1675}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_3128, signal_469}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_94 ( .s (signal_457), .b ({signal_2165, signal_1674}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_3129, signal_471}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_97 ( .s (signal_457), .b ({signal_2168, signal_1673}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_3130, signal_473}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_100 ( .s (signal_457), .b ({signal_2171, signal_1672}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_3131, signal_475}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_103 ( .s (signal_457), .b ({signal_2174, signal_1671}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_3132, signal_477}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_106 ( .s (signal_457), .b ({signal_2177, signal_1670}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_3133, signal_479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_109 ( .s (signal_457), .b ({signal_2180, signal_1669}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_3134, signal_481}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_112 ( .s (signal_457), .b ({signal_2183, signal_1668}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_3135, signal_483}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_115 ( .s (signal_457), .b ({signal_2186, signal_1667}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_3136, signal_485}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_118 ( .s (signal_457), .b ({signal_2189, signal_1666}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_3137, signal_487}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_121 ( .s (signal_457), .b ({signal_2192, signal_1665}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_3138, signal_489}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_124 ( .s (signal_457), .b ({signal_2195, signal_1664}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_3139, signal_491}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_127 ( .s (signal_457), .b ({signal_2198, signal_1663}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_3140, signal_493}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_130 ( .s (signal_457), .b ({signal_2201, signal_1662}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_3141, signal_495}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_133 ( .s (signal_458), .b ({signal_2204, signal_1661}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_3142, signal_497}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_136 ( .s (signal_458), .b ({signal_2207, signal_1660}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_3143, signal_499}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_139 ( .s (signal_458), .b ({signal_2210, signal_1659}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_3144, signal_501}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_142 ( .s (signal_458), .b ({signal_2213, signal_1658}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_3145, signal_503}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_145 ( .s (signal_458), .b ({signal_2216, signal_1657}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_3146, signal_505}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_148 ( .s (signal_458), .b ({signal_2219, signal_1656}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_3147, signal_507}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_151 ( .s (signal_458), .b ({signal_2222, signal_1655}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_3148, signal_509}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_154 ( .s (signal_458), .b ({signal_2225, signal_1654}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_3149, signal_511}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_157 ( .s (signal_458), .b ({signal_3039, signal_1653}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_3150, signal_513}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_160 ( .s (signal_458), .b ({signal_3041, signal_1652}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_3151, signal_515}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_163 ( .s (signal_458), .b ({signal_3043, signal_1651}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_3152, signal_517}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_166 ( .s (signal_458), .b ({signal_3045, signal_1650}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_3153, signal_519}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_169 ( .s (signal_458), .b ({signal_3047, signal_1649}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_3154, signal_521}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_172 ( .s (signal_458), .b ({signal_3049, signal_1648}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_3155, signal_523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_175 ( .s (signal_458), .b ({signal_3051, signal_1647}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_3156, signal_525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_178 ( .s (signal_458), .b ({signal_3053, signal_1646}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_3157, signal_527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_181 ( .s (signal_459), .b ({signal_2228, signal_1645}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_3158, signal_529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_184 ( .s (signal_459), .b ({signal_2231, signal_1644}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_3159, signal_531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_187 ( .s (signal_459), .b ({signal_2234, signal_1643}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_3160, signal_533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_190 ( .s (signal_459), .b ({signal_2237, signal_1642}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_3161, signal_535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_193 ( .s (signal_459), .b ({signal_2240, signal_1641}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_3162, signal_537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_196 ( .s (signal_459), .b ({signal_2243, signal_1640}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_3163, signal_539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_199 ( .s (signal_459), .b ({signal_2246, signal_1639}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_3164, signal_541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_202 ( .s (signal_459), .b ({signal_2249, signal_1638}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_3165, signal_543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_205 ( .s (signal_459), .b ({signal_2252, signal_1637}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_3166, signal_545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_208 ( .s (signal_459), .b ({signal_2255, signal_1636}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_3167, signal_547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_211 ( .s (signal_459), .b ({signal_2258, signal_1635}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_3168, signal_549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_214 ( .s (signal_459), .b ({signal_2261, signal_1634}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_3169, signal_551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_217 ( .s (signal_459), .b ({signal_2264, signal_1633}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_3170, signal_553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_220 ( .s (signal_459), .b ({signal_2267, signal_1632}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_3171, signal_555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_223 ( .s (signal_459), .b ({signal_2270, signal_1631}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_3172, signal_557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_226 ( .s (signal_459), .b ({signal_2273, signal_1630}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_3173, signal_559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_229 ( .s (signal_460), .b ({signal_2276, signal_1629}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_3174, signal_561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_232 ( .s (signal_460), .b ({signal_2279, signal_1628}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_3175, signal_563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_235 ( .s (signal_460), .b ({signal_2282, signal_1627}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_3176, signal_565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_238 ( .s (signal_460), .b ({signal_2285, signal_1626}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_3177, signal_567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_241 ( .s (signal_460), .b ({signal_2288, signal_1625}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_3178, signal_569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_244 ( .s (signal_460), .b ({signal_2291, signal_1624}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_3179, signal_571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_247 ( .s (signal_460), .b ({signal_2294, signal_1623}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_3180, signal_573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_250 ( .s (signal_460), .b ({signal_2297, signal_1622}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_3181, signal_575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_253 ( .s (signal_460), .b ({signal_3055, signal_1621}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_3182, signal_577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_256 ( .s (signal_460), .b ({signal_3057, signal_1620}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_3183, signal_579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_259 ( .s (signal_460), .b ({signal_3059, signal_1619}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_3184, signal_581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_262 ( .s (signal_460), .b ({signal_3061, signal_1618}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_3185, signal_583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_265 ( .s (signal_460), .b ({signal_3063, signal_1617}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_3186, signal_585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_268 ( .s (signal_460), .b ({signal_3065, signal_1616}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_3187, signal_587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_271 ( .s (signal_460), .b ({signal_3067, signal_1615}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_3188, signal_589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_274 ( .s (signal_460), .b ({signal_3069, signal_1614}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_3189, signal_591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_277 ( .s (signal_461), .b ({signal_2300, signal_1613}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_3190, signal_593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_280 ( .s (signal_461), .b ({signal_2303, signal_1612}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_3191, signal_595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_283 ( .s (signal_461), .b ({signal_2306, signal_1611}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_3192, signal_597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_286 ( .s (signal_461), .b ({signal_2309, signal_1610}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_3193, signal_599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_289 ( .s (signal_461), .b ({signal_2312, signal_1609}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_3194, signal_601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_292 ( .s (signal_461), .b ({signal_2315, signal_1608}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_3195, signal_603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_295 ( .s (signal_461), .b ({signal_2318, signal_1607}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_3196, signal_605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_298 ( .s (signal_461), .b ({signal_2321, signal_1606}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_3197, signal_607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_301 ( .s (signal_461), .b ({signal_2324, signal_1605}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_3198, signal_609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_304 ( .s (signal_461), .b ({signal_2327, signal_1604}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_3199, signal_611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_307 ( .s (signal_461), .b ({signal_2330, signal_1603}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_3200, signal_613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_310 ( .s (signal_461), .b ({signal_2333, signal_1602}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_3201, signal_615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_313 ( .s (signal_461), .b ({signal_2336, signal_1601}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_3202, signal_617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_316 ( .s (signal_461), .b ({signal_2339, signal_1600}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_3203, signal_619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_319 ( .s (signal_461), .b ({signal_2342, signal_1599}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_3204, signal_621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_322 ( .s (signal_461), .b ({signal_2345, signal_1598}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_3205, signal_623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_325 ( .s (signal_462), .b ({signal_2348, signal_1597}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_3206, signal_625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_328 ( .s (signal_462), .b ({signal_2351, signal_1596}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_3207, signal_627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_331 ( .s (signal_462), .b ({signal_2354, signal_1595}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_3208, signal_629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_334 ( .s (signal_462), .b ({signal_2357, signal_1594}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_3209, signal_631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_337 ( .s (signal_462), .b ({signal_2360, signal_1593}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_3210, signal_633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_340 ( .s (signal_462), .b ({signal_2363, signal_1592}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_3211, signal_635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_343 ( .s (signal_462), .b ({signal_2366, signal_1591}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_3212, signal_637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_346 ( .s (signal_462), .b ({signal_2369, signal_1590}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_3213, signal_639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_349 ( .s (signal_462), .b ({signal_3071, signal_1589}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_3214, signal_641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_352 ( .s (signal_462), .b ({signal_3073, signal_1588}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_3215, signal_643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_355 ( .s (signal_462), .b ({signal_3075, signal_1587}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_3216, signal_645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_358 ( .s (signal_462), .b ({signal_3077, signal_1586}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_3217, signal_647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_361 ( .s (signal_462), .b ({signal_3079, signal_1585}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_3218, signal_649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_364 ( .s (signal_462), .b ({signal_3081, signal_1584}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_3219, signal_651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_367 ( .s (signal_462), .b ({signal_3083, signal_1583}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_3220, signal_653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_370 ( .s (signal_462), .b ({signal_3085, signal_1582}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_3221, signal_655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_373 ( .s (signal_463), .b ({signal_2372, signal_1581}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_3222, signal_657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_376 ( .s (signal_463), .b ({signal_2375, signal_1580}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_3223, signal_659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_379 ( .s (signal_463), .b ({signal_2378, signal_1579}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_3224, signal_661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_382 ( .s (signal_463), .b ({signal_2381, signal_1578}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_3225, signal_663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_385 ( .s (signal_463), .b ({signal_2384, signal_1577}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_3226, signal_665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_388 ( .s (signal_463), .b ({signal_2387, signal_1576}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_3227, signal_667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_391 ( .s (signal_463), .b ({signal_2390, signal_1575}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_3228, signal_669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_394 ( .s (signal_463), .b ({signal_2393, signal_1574}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_3229, signal_671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_397 ( .s (signal_463), .b ({signal_2396, signal_1573}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_3230, signal_673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_400 ( .s (signal_463), .b ({signal_2399, signal_1572}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_3231, signal_675}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_403 ( .s (signal_463), .b ({signal_2402, signal_1571}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_3232, signal_677}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_406 ( .s (signal_463), .b ({signal_2405, signal_1570}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_3233, signal_679}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_409 ( .s (signal_463), .b ({signal_2408, signal_1569}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_3234, signal_681}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_412 ( .s (signal_463), .b ({signal_2411, signal_1568}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_3235, signal_683}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_415 ( .s (signal_463), .b ({signal_2414, signal_1567}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_3236, signal_685}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_418 ( .s (signal_463), .b ({signal_2417, signal_1566}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_3237, signal_687}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_421 ( .s (signal_464), .b ({signal_2420, signal_1565}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_3238, signal_689}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_424 ( .s (signal_464), .b ({signal_2423, signal_1564}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_3239, signal_691}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_427 ( .s (signal_464), .b ({signal_2426, signal_1563}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_3240, signal_693}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_430 ( .s (signal_464), .b ({signal_2429, signal_1562}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_3241, signal_695}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_433 ( .s (signal_464), .b ({signal_2432, signal_1561}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_3242, signal_697}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_436 ( .s (signal_464), .b ({signal_2435, signal_1560}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_3243, signal_699}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_439 ( .s (signal_464), .b ({signal_2438, signal_1559}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_3244, signal_701}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_442 ( .s (signal_464), .b ({signal_2441, signal_1558}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_3245, signal_703}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_469 ( .s (signal_445), .b ({plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_2156, signal_1677}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_470 ( .s (signal_445), .b ({plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_2159, signal_1676}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_471 ( .s (signal_445), .b ({plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_2162, signal_1675}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_472 ( .s (signal_445), .b ({plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_2165, signal_1674}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_473 ( .s (signal_445), .b ({plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_2168, signal_1673}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_474 ( .s (signal_445), .b ({plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_2171, signal_1672}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_475 ( .s (signal_445), .b ({plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_2174, signal_1671}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_476 ( .s (signal_445), .b ({plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_2177, signal_1670}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_477 ( .s (signal_445), .b ({plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_2180, signal_1669}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_478 ( .s (signal_445), .b ({plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_2183, signal_1668}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_479 ( .s (signal_445), .b ({plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_2186, signal_1667}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_480 ( .s (signal_445), .b ({plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_2189, signal_1666}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_481 ( .s (signal_445), .b ({plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_2192, signal_1665}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_482 ( .s (signal_445), .b ({plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_2195, signal_1664}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_483 ( .s (signal_445), .b ({plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_2198, signal_1663}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_484 ( .s (signal_445), .b ({plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_2201, signal_1662}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_485 ( .s (signal_446), .b ({plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_2204, signal_1661}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_486 ( .s (signal_446), .b ({plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_2207, signal_1660}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_487 ( .s (signal_446), .b ({plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_2210, signal_1659}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_488 ( .s (signal_446), .b ({plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_2213, signal_1658}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_489 ( .s (signal_446), .b ({plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_2216, signal_1657}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_490 ( .s (signal_446), .b ({plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_2219, signal_1656}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_491 ( .s (signal_446), .b ({plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_2222, signal_1655}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_492 ( .s (signal_446), .b ({plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_2225, signal_1654}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_493 ( .s (signal_454), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_2870, signal_1429}), .c ({signal_3006, signal_1549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_494 ( .s (signal_454), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_2871, signal_1428}), .c ({signal_3007, signal_1548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_495 ( .s (signal_454), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_2872, signal_1427}), .c ({signal_3008, signal_1547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_496 ( .s (signal_454), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_2873, signal_1426}), .c ({signal_3009, signal_1546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_497 ( .s (signal_454), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_2874, signal_1425}), .c ({signal_3010, signal_1545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_498 ( .s (signal_454), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_2875, signal_1424}), .c ({signal_3011, signal_1544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_499 ( .s (signal_454), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_2876, signal_1423}), .c ({signal_3012, signal_1543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_500 ( .s (signal_454), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_2877, signal_1422}), .c ({signal_3013, signal_1542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_501 ( .s (signal_446), .b ({plaintext_s1[96], plaintext_s0[96]}), .a ({signal_3006, signal_1549}), .c ({signal_3039, signal_1653}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_502 ( .s (signal_446), .b ({plaintext_s1[97], plaintext_s0[97]}), .a ({signal_3007, signal_1548}), .c ({signal_3041, signal_1652}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_503 ( .s (signal_446), .b ({plaintext_s1[98], plaintext_s0[98]}), .a ({signal_3008, signal_1547}), .c ({signal_3043, signal_1651}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_504 ( .s (signal_446), .b ({plaintext_s1[99], plaintext_s0[99]}), .a ({signal_3009, signal_1546}), .c ({signal_3045, signal_1650}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_505 ( .s (signal_446), .b ({plaintext_s1[100], plaintext_s0[100]}), .a ({signal_3010, signal_1545}), .c ({signal_3047, signal_1649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_506 ( .s (signal_446), .b ({plaintext_s1[101], plaintext_s0[101]}), .a ({signal_3011, signal_1544}), .c ({signal_3049, signal_1648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_507 ( .s (signal_446), .b ({plaintext_s1[102], plaintext_s0[102]}), .a ({signal_3012, signal_1543}), .c ({signal_3051, signal_1647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_508 ( .s (signal_446), .b ({plaintext_s1[103], plaintext_s0[103]}), .a ({signal_3013, signal_1542}), .c ({signal_3053, signal_1646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_509 ( .s (signal_447), .b ({plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_2228, signal_1645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_510 ( .s (signal_447), .b ({plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_2231, signal_1644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_511 ( .s (signal_447), .b ({plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_2234, signal_1643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_512 ( .s (signal_447), .b ({plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_2237, signal_1642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_513 ( .s (signal_447), .b ({plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_2240, signal_1641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_514 ( .s (signal_447), .b ({plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_2243, signal_1640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_515 ( .s (signal_447), .b ({plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_2246, signal_1639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_516 ( .s (signal_447), .b ({plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_2249, signal_1638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_517 ( .s (signal_447), .b ({plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_2252, signal_1637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_518 ( .s (signal_447), .b ({plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_2255, signal_1636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_519 ( .s (signal_447), .b ({plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_2258, signal_1635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_520 ( .s (signal_447), .b ({plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_2261, signal_1634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_521 ( .s (signal_447), .b ({plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_2264, signal_1633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_522 ( .s (signal_447), .b ({plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_2267, signal_1632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_523 ( .s (signal_447), .b ({plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_2270, signal_1631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_524 ( .s (signal_447), .b ({plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_2273, signal_1630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_525 ( .s (signal_448), .b ({plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_2276, signal_1629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_526 ( .s (signal_448), .b ({plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_2279, signal_1628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_527 ( .s (signal_448), .b ({plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_2282, signal_1627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_528 ( .s (signal_448), .b ({plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_2285, signal_1626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_529 ( .s (signal_448), .b ({plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_2288, signal_1625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_530 ( .s (signal_448), .b ({plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_2291, signal_1624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_531 ( .s (signal_448), .b ({plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_2294, signal_1623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_532 ( .s (signal_448), .b ({plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_2297, signal_1622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_533 ( .s (signal_454), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_2862, signal_1437}), .c ({signal_3014, signal_1541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_534 ( .s (signal_454), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_2863, signal_1436}), .c ({signal_3015, signal_1540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_535 ( .s (signal_454), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_2864, signal_1435}), .c ({signal_3016, signal_1539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_536 ( .s (signal_454), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_2865, signal_1434}), .c ({signal_3017, signal_1538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_537 ( .s (signal_454), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_2866, signal_1433}), .c ({signal_3018, signal_1537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_538 ( .s (signal_454), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_2867, signal_1432}), .c ({signal_3019, signal_1536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_539 ( .s (signal_454), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_2868, signal_1431}), .c ({signal_3020, signal_1535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_540 ( .s (signal_454), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_2869, signal_1430}), .c ({signal_3021, signal_1534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_541 ( .s (signal_448), .b ({plaintext_s1[64], plaintext_s0[64]}), .a ({signal_3014, signal_1541}), .c ({signal_3055, signal_1621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_542 ( .s (signal_448), .b ({plaintext_s1[65], plaintext_s0[65]}), .a ({signal_3015, signal_1540}), .c ({signal_3057, signal_1620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_543 ( .s (signal_448), .b ({plaintext_s1[66], plaintext_s0[66]}), .a ({signal_3016, signal_1539}), .c ({signal_3059, signal_1619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_544 ( .s (signal_448), .b ({plaintext_s1[67], plaintext_s0[67]}), .a ({signal_3017, signal_1538}), .c ({signal_3061, signal_1618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_545 ( .s (signal_448), .b ({plaintext_s1[68], plaintext_s0[68]}), .a ({signal_3018, signal_1537}), .c ({signal_3063, signal_1617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_546 ( .s (signal_448), .b ({plaintext_s1[69], plaintext_s0[69]}), .a ({signal_3019, signal_1536}), .c ({signal_3065, signal_1616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_547 ( .s (signal_448), .b ({plaintext_s1[70], plaintext_s0[70]}), .a ({signal_3020, signal_1535}), .c ({signal_3067, signal_1615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_548 ( .s (signal_448), .b ({plaintext_s1[71], plaintext_s0[71]}), .a ({signal_3021, signal_1534}), .c ({signal_3069, signal_1614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_549 ( .s (signal_449), .b ({plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_2300, signal_1613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_550 ( .s (signal_449), .b ({plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_2303, signal_1612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_551 ( .s (signal_449), .b ({plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_2306, signal_1611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_552 ( .s (signal_449), .b ({plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_2309, signal_1610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_553 ( .s (signal_449), .b ({plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_2312, signal_1609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_554 ( .s (signal_449), .b ({plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_2315, signal_1608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_555 ( .s (signal_449), .b ({plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_2318, signal_1607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_556 ( .s (signal_449), .b ({plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_2321, signal_1606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_557 ( .s (signal_449), .b ({plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_2324, signal_1605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_558 ( .s (signal_449), .b ({plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_2327, signal_1604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_559 ( .s (signal_449), .b ({plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_2330, signal_1603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_560 ( .s (signal_449), .b ({plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_2333, signal_1602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_561 ( .s (signal_449), .b ({plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_2336, signal_1601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_562 ( .s (signal_449), .b ({plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_2339, signal_1600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_563 ( .s (signal_449), .b ({plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_2342, signal_1599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_564 ( .s (signal_449), .b ({plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_2345, signal_1598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_565 ( .s (signal_450), .b ({plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_2348, signal_1597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_566 ( .s (signal_450), .b ({plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_2351, signal_1596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_567 ( .s (signal_450), .b ({plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_2354, signal_1595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_568 ( .s (signal_450), .b ({plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_2357, signal_1594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_569 ( .s (signal_450), .b ({plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_2360, signal_1593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_570 ( .s (signal_450), .b ({plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_2363, signal_1592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_571 ( .s (signal_450), .b ({plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_2366, signal_1591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_572 ( .s (signal_450), .b ({plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_2369, signal_1590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_573 ( .s (signal_455), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_2854, signal_1445}), .c ({signal_3022, signal_1533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_574 ( .s (signal_455), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_2855, signal_1444}), .c ({signal_3023, signal_1532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_575 ( .s (signal_455), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_2856, signal_1443}), .c ({signal_3024, signal_1531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_576 ( .s (signal_455), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_2857, signal_1442}), .c ({signal_3025, signal_1530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_577 ( .s (signal_455), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_2858, signal_1441}), .c ({signal_3026, signal_1529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_578 ( .s (signal_455), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_2859, signal_1440}), .c ({signal_3027, signal_1528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_579 ( .s (signal_455), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_2860, signal_1439}), .c ({signal_3028, signal_1527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_580 ( .s (signal_455), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_2861, signal_1438}), .c ({signal_3029, signal_1526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_581 ( .s (signal_450), .b ({plaintext_s1[32], plaintext_s0[32]}), .a ({signal_3022, signal_1533}), .c ({signal_3071, signal_1589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_582 ( .s (signal_450), .b ({plaintext_s1[33], plaintext_s0[33]}), .a ({signal_3023, signal_1532}), .c ({signal_3073, signal_1588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_583 ( .s (signal_450), .b ({plaintext_s1[34], plaintext_s0[34]}), .a ({signal_3024, signal_1531}), .c ({signal_3075, signal_1587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_584 ( .s (signal_450), .b ({plaintext_s1[35], plaintext_s0[35]}), .a ({signal_3025, signal_1530}), .c ({signal_3077, signal_1586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_585 ( .s (signal_450), .b ({plaintext_s1[36], plaintext_s0[36]}), .a ({signal_3026, signal_1529}), .c ({signal_3079, signal_1585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_586 ( .s (signal_450), .b ({plaintext_s1[37], plaintext_s0[37]}), .a ({signal_3027, signal_1528}), .c ({signal_3081, signal_1584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_587 ( .s (signal_450), .b ({plaintext_s1[38], plaintext_s0[38]}), .a ({signal_3028, signal_1527}), .c ({signal_3083, signal_1583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_588 ( .s (signal_450), .b ({plaintext_s1[39], plaintext_s0[39]}), .a ({signal_3029, signal_1526}), .c ({signal_3085, signal_1582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_589 ( .s (signal_451), .b ({plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_2372, signal_1581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_590 ( .s (signal_451), .b ({plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_2375, signal_1580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_591 ( .s (signal_451), .b ({plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_2378, signal_1579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_592 ( .s (signal_451), .b ({plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_2381, signal_1578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_593 ( .s (signal_451), .b ({plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_2384, signal_1577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_594 ( .s (signal_451), .b ({plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_2387, signal_1576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_595 ( .s (signal_451), .b ({plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_2390, signal_1575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_596 ( .s (signal_451), .b ({plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_2393, signal_1574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_597 ( .s (signal_451), .b ({plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_2396, signal_1573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_598 ( .s (signal_451), .b ({plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_2399, signal_1572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_599 ( .s (signal_451), .b ({plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({signal_2402, signal_1571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_600 ( .s (signal_451), .b ({plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({signal_2405, signal_1570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_601 ( .s (signal_451), .b ({plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_2408, signal_1569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_602 ( .s (signal_451), .b ({plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_2411, signal_1568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_603 ( .s (signal_451), .b ({plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_2414, signal_1567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_604 ( .s (signal_451), .b ({plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_2417, signal_1566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_605 ( .s (signal_452), .b ({plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_2420, signal_1565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_606 ( .s (signal_452), .b ({plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_2423, signal_1564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_607 ( .s (signal_452), .b ({plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_2426, signal_1563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_608 ( .s (signal_452), .b ({plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_2429, signal_1562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_609 ( .s (signal_452), .b ({plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_2432, signal_1561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_610 ( .s (signal_452), .b ({plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_2435, signal_1560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_611 ( .s (signal_452), .b ({plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_2438, signal_1559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_612 ( .s (signal_452), .b ({plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_2441, signal_1558}) ) ;
    INV_X1 cell_629 ( .A (signal_399), .ZN (signal_721) ) ;
    INV_X1 cell_630 ( .A (signal_721), .ZN (signal_722) ) ;
    INV_X1 cell_631 ( .A (signal_721), .ZN (signal_723) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_632 ( .s (signal_723), .b ({signal_2825, signal_1485}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2850, signal_1453}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_633 ( .s (signal_722), .b ({signal_2849, signal_1484}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2851, signal_1452}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_634 ( .s (signal_399), .b ({signal_2823, signal_1483}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2834, signal_1451}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_635 ( .s (signal_399), .b ({signal_2848, signal_1482}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2852, signal_1450}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_636 ( .s (signal_399), .b ({signal_2847, signal_1481}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2853, signal_1449}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_637 ( .s (signal_399), .b ({signal_2820, signal_1480}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2835, signal_1448}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_638 ( .s (signal_399), .b ({signal_2819, signal_1479}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2836, signal_1447}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_639 ( .s (signal_399), .b ({signal_2818, signal_1478}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2837, signal_1446}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_640 ( .s (signal_722), .b ({signal_2817, signal_1477}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2854, signal_1445}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_641 ( .s (signal_722), .b ({signal_2846, signal_1476}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2855, signal_1444}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_642 ( .s (signal_722), .b ({signal_2815, signal_1475}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2856, signal_1443}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_643 ( .s (signal_722), .b ({signal_2845, signal_1474}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2857, signal_1442}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_644 ( .s (signal_722), .b ({signal_2844, signal_1473}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2858, signal_1441}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_645 ( .s (signal_722), .b ({signal_2812, signal_1472}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2859, signal_1440}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_646 ( .s (signal_722), .b ({signal_2811, signal_1471}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2860, signal_1439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_647 ( .s (signal_722), .b ({signal_2810, signal_1470}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2861, signal_1438}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_648 ( .s (signal_722), .b ({signal_2809, signal_1469}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2862, signal_1437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_649 ( .s (signal_722), .b ({signal_2843, signal_1468}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2863, signal_1436}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_650 ( .s (signal_722), .b ({signal_2807, signal_1467}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2864, signal_1435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_651 ( .s (signal_722), .b ({signal_2842, signal_1466}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2865, signal_1434}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_652 ( .s (signal_723), .b ({signal_2841, signal_1465}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2866, signal_1433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_653 ( .s (signal_723), .b ({signal_2804, signal_1464}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2867, signal_1432}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_654 ( .s (signal_723), .b ({signal_2803, signal_1463}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2868, signal_1431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_655 ( .s (signal_723), .b ({signal_2802, signal_1462}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2869, signal_1430}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_656 ( .s (signal_723), .b ({signal_2801, signal_1461}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2870, signal_1429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_657 ( .s (signal_723), .b ({signal_2840, signal_1460}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2871, signal_1428}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_658 ( .s (signal_723), .b ({signal_2799, signal_1459}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2872, signal_1427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_659 ( .s (signal_723), .b ({signal_2839, signal_1458}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2873, signal_1426}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_660 ( .s (signal_723), .b ({signal_2838, signal_1457}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2874, signal_1425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_661 ( .s (signal_723), .b ({signal_2796, signal_1456}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2875, signal_1424}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_662 ( .s (signal_723), .b ({signal_2795, signal_1455}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2876, signal_1423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_663 ( .s (signal_723), .b ({signal_2794, signal_1454}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2877, signal_1422}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_664 ( .a ({signal_2006, signal_765}), .b ({signal_2004, signal_1486}), .c ({signal_2007, signal_1686}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_665 ( .a ({signal_2008, signal_764}), .b ({signal_2001, signal_1487}), .c ({signal_2009, signal_1687}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_666 ( .a ({signal_2010, signal_763}), .b ({signal_1998, signal_1488}), .c ({signal_2011, signal_1688}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_667 ( .a ({signal_2012, signal_762}), .b ({signal_1995, signal_1489}), .c ({signal_2013, signal_1689}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_668 ( .a ({signal_2014, signal_761}), .b ({signal_1992, signal_1490}), .c ({signal_2015, signal_1690}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_669 ( .a ({signal_2016, signal_760}), .b ({signal_1989, signal_1491}), .c ({signal_2017, signal_1691}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_670 ( .a ({signal_2018, signal_759}), .b ({signal_1986, signal_1492}), .c ({signal_2019, signal_1692}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_671 ( .a ({signal_2020, signal_758}), .b ({signal_1983, signal_1493}), .c ({signal_2021, signal_1693}) ) ;
    INV_X1 cell_688 ( .A (signal_732), .ZN (signal_733) ) ;
    INV_X1 cell_689 ( .A (signal_732), .ZN (signal_734) ) ;
    INV_X1 cell_690 ( .A (signal_732), .ZN (signal_735) ) ;
    INV_X1 cell_691 ( .A (signal_732), .ZN (signal_736) ) ;
    INV_X1 cell_692 ( .A (signal_732), .ZN (signal_737) ) ;
    INV_X1 cell_693 ( .A (signal_732), .ZN (signal_738) ) ;
    INV_X1 cell_694 ( .A (signal_732), .ZN (signal_739) ) ;
    INV_X1 cell_695 ( .A (signal_732), .ZN (signal_740) ) ;
    INV_X1 cell_696 ( .A (signal_393), .ZN (signal_732) ) ;
    INV_X1 cell_697 ( .A (signal_741), .ZN (signal_748) ) ;
    INV_X1 cell_698 ( .A (signal_750), .ZN (signal_756) ) ;
    INV_X1 cell_699 ( .A (signal_741), .ZN (signal_742) ) ;
    INV_X1 cell_700 ( .A (signal_750), .ZN (signal_751) ) ;
    INV_X1 cell_701 ( .A (signal_741), .ZN (signal_743) ) ;
    INV_X1 cell_702 ( .A (signal_750), .ZN (signal_752) ) ;
    INV_X1 cell_703 ( .A (signal_741), .ZN (signal_744) ) ;
    INV_X1 cell_704 ( .A (signal_750), .ZN (signal_753) ) ;
    INV_X1 cell_705 ( .A (signal_741), .ZN (signal_747) ) ;
    INV_X1 cell_706 ( .A (signal_750), .ZN (signal_755) ) ;
    INV_X1 cell_707 ( .A (signal_741), .ZN (signal_746) ) ;
    INV_X1 cell_708 ( .A (signal_750), .ZN (signal_754) ) ;
    INV_X1 cell_709 ( .A (signal_741), .ZN (signal_749) ) ;
    INV_X1 cell_710 ( .A (signal_750), .ZN (signal_757) ) ;
    INV_X1 cell_711 ( .A (signal_741), .ZN (signal_745) ) ;
    INV_X1 cell_712 ( .A (signal_394), .ZN (signal_741) ) ;
    INV_X1 cell_713 ( .A (signal_404), .ZN (signal_750) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_714 ( .s (signal_751), .b ({signal_1983, signal_1493}), .a ({signal_3294, signal_767}), .c ({signal_3406, signal_766}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_715 ( .s (signal_742), .b ({signal_3271, signal_1933}), .a ({signal_2491, signal_1877}), .c ({signal_3294, signal_767}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_718 ( .s (signal_751), .b ({signal_1986, signal_1492}), .a ({signal_3295, signal_770}), .c ({signal_3407, signal_769}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_719 ( .s (signal_742), .b ({signal_3273, signal_1932}), .a ({signal_2494, signal_1876}), .c ({signal_3295, signal_770}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_722 ( .s (signal_751), .b ({signal_1989, signal_1491}), .a ({signal_3296, signal_773}), .c ({signal_3408, signal_772}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_723 ( .s (signal_742), .b ({signal_3275, signal_1931}), .a ({signal_2497, signal_1875}), .c ({signal_3296, signal_773}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_726 ( .s (signal_751), .b ({signal_1992, signal_1490}), .a ({signal_3297, signal_776}), .c ({signal_3409, signal_775}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_727 ( .s (signal_742), .b ({signal_3277, signal_1930}), .a ({signal_2500, signal_1874}), .c ({signal_3297, signal_776}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_730 ( .s (signal_751), .b ({signal_1995, signal_1489}), .a ({signal_3298, signal_779}), .c ({signal_3410, signal_778}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_731 ( .s (signal_742), .b ({signal_3279, signal_1929}), .a ({signal_2503, signal_1873}), .c ({signal_3298, signal_779}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_734 ( .s (signal_751), .b ({signal_1998, signal_1488}), .a ({signal_3299, signal_782}), .c ({signal_3411, signal_781}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_735 ( .s (signal_742), .b ({signal_3281, signal_1928}), .a ({signal_2506, signal_1872}), .c ({signal_3299, signal_782}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_738 ( .s (signal_751), .b ({signal_2001, signal_1487}), .a ({signal_3300, signal_785}), .c ({signal_3412, signal_784}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_739 ( .s (signal_742), .b ({signal_3283, signal_1927}), .a ({signal_2509, signal_1871}), .c ({signal_3300, signal_785}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_742 ( .s (signal_751), .b ({signal_2004, signal_1486}), .a ({signal_3301, signal_788}), .c ({signal_3413, signal_787}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_743 ( .s (signal_742), .b ({signal_3285, signal_1926}), .a ({signal_2512, signal_1870}), .c ({signal_3301, signal_788}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_746 ( .s (signal_751), .b ({signal_2020, signal_758}), .a ({signal_2878, signal_791}), .c ({signal_3302, signal_790}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_747 ( .s (signal_742), .b ({signal_2444, signal_1925}), .a ({signal_2515, signal_1861}), .c ({signal_2878, signal_791}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_750 ( .s (signal_751), .b ({signal_2018, signal_759}), .a ({signal_2879, signal_794}), .c ({signal_3303, signal_793}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_751 ( .s (signal_742), .b ({signal_2447, signal_1924}), .a ({signal_2518, signal_1860}), .c ({signal_2879, signal_794}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_754 ( .s (signal_751), .b ({signal_2016, signal_760}), .a ({signal_2880, signal_797}), .c ({signal_3304, signal_796}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_755 ( .s (signal_742), .b ({signal_2450, signal_1923}), .a ({signal_2521, signal_1859}), .c ({signal_2880, signal_797}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_758 ( .s (signal_751), .b ({signal_2014, signal_761}), .a ({signal_2881, signal_800}), .c ({signal_3305, signal_799}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_759 ( .s (signal_742), .b ({signal_2453, signal_1922}), .a ({signal_2524, signal_1858}), .c ({signal_2881, signal_800}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_762 ( .s (signal_751), .b ({signal_2012, signal_762}), .a ({signal_2882, signal_803}), .c ({signal_3306, signal_802}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_763 ( .s (signal_742), .b ({signal_2456, signal_1921}), .a ({signal_2527, signal_1857}), .c ({signal_2882, signal_803}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_766 ( .s (signal_751), .b ({signal_2010, signal_763}), .a ({signal_2883, signal_806}), .c ({signal_3307, signal_805}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_767 ( .s (signal_742), .b ({signal_2459, signal_1920}), .a ({signal_2530, signal_1856}), .c ({signal_2883, signal_806}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_770 ( .s (signal_751), .b ({signal_2008, signal_764}), .a ({signal_2884, signal_809}), .c ({signal_3308, signal_808}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_771 ( .s (signal_742), .b ({signal_2462, signal_1919}), .a ({signal_2533, signal_1855}), .c ({signal_2884, signal_809}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_774 ( .s (signal_751), .b ({signal_2006, signal_765}), .a ({signal_2885, signal_812}), .c ({signal_3309, signal_811}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_775 ( .s (signal_742), .b ({signal_2465, signal_1918}), .a ({signal_2536, signal_1854}), .c ({signal_2885, signal_812}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_778 ( .s (signal_752), .b ({signal_2443, signal_1909}), .a ({signal_2886, signal_815}), .c ({signal_3310, signal_814}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_779 ( .s (signal_743), .b ({signal_2468, signal_1917}), .a ({signal_2539, signal_1845}), .c ({signal_2886, signal_815}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_782 ( .s (signal_752), .b ({signal_2446, signal_1908}), .a ({signal_2887, signal_818}), .c ({signal_3311, signal_817}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_783 ( .s (signal_743), .b ({signal_2471, signal_1916}), .a ({signal_2542, signal_1844}), .c ({signal_2887, signal_818}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_786 ( .s (signal_752), .b ({signal_2449, signal_1907}), .a ({signal_2888, signal_821}), .c ({signal_3312, signal_820}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_787 ( .s (signal_743), .b ({signal_2474, signal_1915}), .a ({signal_2545, signal_1843}), .c ({signal_2888, signal_821}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_790 ( .s (signal_752), .b ({signal_2452, signal_1906}), .a ({signal_2889, signal_824}), .c ({signal_3313, signal_823}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_791 ( .s (signal_743), .b ({signal_2477, signal_1914}), .a ({signal_2548, signal_1842}), .c ({signal_2889, signal_824}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_794 ( .s (signal_752), .b ({signal_2455, signal_1905}), .a ({signal_2890, signal_827}), .c ({signal_3314, signal_826}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_795 ( .s (signal_743), .b ({signal_2480, signal_1913}), .a ({signal_2551, signal_1841}), .c ({signal_2890, signal_827}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_798 ( .s (signal_752), .b ({signal_2458, signal_1904}), .a ({signal_2891, signal_830}), .c ({signal_3315, signal_829}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_799 ( .s (signal_743), .b ({signal_2483, signal_1912}), .a ({signal_2554, signal_1840}), .c ({signal_2891, signal_830}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_802 ( .s (signal_752), .b ({signal_2461, signal_1903}), .a ({signal_2892, signal_833}), .c ({signal_3316, signal_832}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_803 ( .s (signal_743), .b ({signal_2486, signal_1911}), .a ({signal_2557, signal_1839}), .c ({signal_2892, signal_833}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_806 ( .s (signal_752), .b ({signal_2464, signal_1902}), .a ({signal_2893, signal_836}), .c ({signal_3317, signal_835}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_807 ( .s (signal_743), .b ({signal_2489, signal_1910}), .a ({signal_2560, signal_1838}), .c ({signal_2893, signal_836}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_810 ( .s (signal_752), .b ({signal_2467, signal_1893}), .a ({signal_2894, signal_839}), .c ({signal_3318, signal_838}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_811 ( .s (signal_743), .b ({signal_2492, signal_1901}), .a ({signal_2563, signal_1509}), .c ({signal_2894, signal_839}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_814 ( .s (signal_752), .b ({signal_2470, signal_1892}), .a ({signal_2895, signal_842}), .c ({signal_3319, signal_841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_815 ( .s (signal_743), .b ({signal_2495, signal_1900}), .a ({signal_2566, signal_1508}), .c ({signal_2895, signal_842}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_818 ( .s (signal_752), .b ({signal_2473, signal_1891}), .a ({signal_2896, signal_845}), .c ({signal_3320, signal_844}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_819 ( .s (signal_743), .b ({signal_2498, signal_1899}), .a ({signal_2569, signal_1507}), .c ({signal_2896, signal_845}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_822 ( .s (signal_752), .b ({signal_2476, signal_1890}), .a ({signal_2897, signal_848}), .c ({signal_3321, signal_847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_823 ( .s (signal_743), .b ({signal_2501, signal_1898}), .a ({signal_2572, signal_1506}), .c ({signal_2897, signal_848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_826 ( .s (signal_752), .b ({signal_2479, signal_1889}), .a ({signal_2898, signal_851}), .c ({signal_3322, signal_850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_827 ( .s (signal_743), .b ({signal_2504, signal_1897}), .a ({signal_2575, signal_1505}), .c ({signal_2898, signal_851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_830 ( .s (signal_752), .b ({signal_2482, signal_1888}), .a ({signal_2899, signal_854}), .c ({signal_3323, signal_853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_831 ( .s (signal_743), .b ({signal_2507, signal_1896}), .a ({signal_2578, signal_1504}), .c ({signal_2899, signal_854}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_834 ( .s (signal_752), .b ({signal_2485, signal_1887}), .a ({signal_2900, signal_857}), .c ({signal_3324, signal_856}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_835 ( .s (signal_743), .b ({signal_2510, signal_1895}), .a ({signal_2581, signal_1503}), .c ({signal_2900, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_838 ( .s (signal_752), .b ({signal_2488, signal_1886}), .a ({signal_2901, signal_860}), .c ({signal_3325, signal_859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_839 ( .s (signal_743), .b ({signal_2513, signal_1894}), .a ({signal_2584, signal_1502}), .c ({signal_2901, signal_860}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_842 ( .s (signal_753), .b ({signal_2491, signal_1877}), .a ({signal_2902, signal_863}), .c ({signal_3326, signal_862}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_843 ( .s (signal_744), .b ({signal_2516, signal_1885}), .a ({signal_2587, signal_1821}), .c ({signal_2902, signal_863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_846 ( .s (signal_753), .b ({signal_2494, signal_1876}), .a ({signal_2903, signal_866}), .c ({signal_3327, signal_865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_847 ( .s (signal_744), .b ({signal_2519, signal_1884}), .a ({signal_2590, signal_1820}), .c ({signal_2903, signal_866}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_850 ( .s (signal_753), .b ({signal_2497, signal_1875}), .a ({signal_2904, signal_869}), .c ({signal_3328, signal_868}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_851 ( .s (signal_744), .b ({signal_2522, signal_1883}), .a ({signal_2593, signal_1819}), .c ({signal_2904, signal_869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_854 ( .s (signal_753), .b ({signal_2500, signal_1874}), .a ({signal_2905, signal_872}), .c ({signal_3329, signal_871}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_855 ( .s (signal_744), .b ({signal_2525, signal_1882}), .a ({signal_2596, signal_1818}), .c ({signal_2905, signal_872}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_858 ( .s (signal_753), .b ({signal_2503, signal_1873}), .a ({signal_2906, signal_875}), .c ({signal_3330, signal_874}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_859 ( .s (signal_744), .b ({signal_2528, signal_1881}), .a ({signal_2599, signal_1817}), .c ({signal_2906, signal_875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_862 ( .s (signal_753), .b ({signal_2506, signal_1872}), .a ({signal_2907, signal_878}), .c ({signal_3331, signal_877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_863 ( .s (signal_744), .b ({signal_2531, signal_1880}), .a ({signal_2602, signal_1816}), .c ({signal_2907, signal_878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_866 ( .s (signal_753), .b ({signal_2509, signal_1871}), .a ({signal_2908, signal_881}), .c ({signal_3332, signal_880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_867 ( .s (signal_744), .b ({signal_2534, signal_1879}), .a ({signal_2605, signal_1815}), .c ({signal_2908, signal_881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_870 ( .s (signal_753), .b ({signal_2512, signal_1870}), .a ({signal_2909, signal_884}), .c ({signal_3333, signal_883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_871 ( .s (signal_744), .b ({signal_2537, signal_1878}), .a ({signal_2608, signal_1814}), .c ({signal_2909, signal_884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_874 ( .s (signal_753), .b ({signal_2515, signal_1861}), .a ({signal_2910, signal_887}), .c ({signal_3334, signal_886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_875 ( .s (signal_744), .b ({signal_2540, signal_1869}), .a ({signal_2611, signal_1805}), .c ({signal_2910, signal_887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_878 ( .s (signal_753), .b ({signal_2518, signal_1860}), .a ({signal_2911, signal_890}), .c ({signal_3335, signal_889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_879 ( .s (signal_744), .b ({signal_2543, signal_1868}), .a ({signal_2614, signal_1804}), .c ({signal_2911, signal_890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_882 ( .s (signal_753), .b ({signal_2521, signal_1859}), .a ({signal_2912, signal_893}), .c ({signal_3336, signal_892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_883 ( .s (signal_744), .b ({signal_2546, signal_1867}), .a ({signal_2617, signal_1803}), .c ({signal_2912, signal_893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_886 ( .s (signal_753), .b ({signal_2524, signal_1858}), .a ({signal_2913, signal_896}), .c ({signal_3337, signal_895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_887 ( .s (signal_744), .b ({signal_2549, signal_1866}), .a ({signal_2620, signal_1802}), .c ({signal_2913, signal_896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_890 ( .s (signal_753), .b ({signal_2527, signal_1857}), .a ({signal_2914, signal_899}), .c ({signal_3338, signal_898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_891 ( .s (signal_744), .b ({signal_2552, signal_1865}), .a ({signal_2623, signal_1801}), .c ({signal_2914, signal_899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_894 ( .s (signal_753), .b ({signal_2530, signal_1856}), .a ({signal_2915, signal_902}), .c ({signal_3339, signal_901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_895 ( .s (signal_744), .b ({signal_2555, signal_1864}), .a ({signal_2626, signal_1800}), .c ({signal_2915, signal_902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_898 ( .s (signal_753), .b ({signal_2533, signal_1855}), .a ({signal_2916, signal_905}), .c ({signal_3340, signal_904}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_899 ( .s (signal_744), .b ({signal_2558, signal_1863}), .a ({signal_2629, signal_1799}), .c ({signal_2916, signal_905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_902 ( .s (signal_753), .b ({signal_2536, signal_1854}), .a ({signal_2917, signal_908}), .c ({signal_3341, signal_907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_903 ( .s (signal_744), .b ({signal_2561, signal_1862}), .a ({signal_2632, signal_1798}), .c ({signal_2917, signal_908}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_906 ( .s (signal_404), .b ({signal_2539, signal_1845}), .a ({signal_2918, signal_911}), .c ({signal_3102, signal_910}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_907 ( .s (signal_745), .b ({signal_2564, signal_1853}), .a ({signal_2635, signal_1789}), .c ({signal_2918, signal_911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_910 ( .s (signal_404), .b ({signal_2542, signal_1844}), .a ({signal_2919, signal_914}), .c ({signal_3103, signal_913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_911 ( .s (signal_745), .b ({signal_2567, signal_1852}), .a ({signal_2638, signal_1788}), .c ({signal_2919, signal_914}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_914 ( .s (signal_404), .b ({signal_2545, signal_1843}), .a ({signal_2920, signal_917}), .c ({signal_3104, signal_916}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_915 ( .s (signal_745), .b ({signal_2570, signal_1851}), .a ({signal_2641, signal_1787}), .c ({signal_2920, signal_917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_918 ( .s (signal_404), .b ({signal_2548, signal_1842}), .a ({signal_2921, signal_920}), .c ({signal_3105, signal_919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_919 ( .s (signal_745), .b ({signal_2573, signal_1850}), .a ({signal_2644, signal_1786}), .c ({signal_2921, signal_920}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_922 ( .s (signal_404), .b ({signal_2551, signal_1841}), .a ({signal_2922, signal_923}), .c ({signal_3106, signal_922}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_923 ( .s (signal_745), .b ({signal_2576, signal_1849}), .a ({signal_2647, signal_1785}), .c ({signal_2922, signal_923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_926 ( .s (signal_404), .b ({signal_2554, signal_1840}), .a ({signal_2923, signal_926}), .c ({signal_3107, signal_925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_927 ( .s (signal_745), .b ({signal_2579, signal_1848}), .a ({signal_2650, signal_1784}), .c ({signal_2923, signal_926}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_930 ( .s (signal_404), .b ({signal_2557, signal_1839}), .a ({signal_2924, signal_929}), .c ({signal_3108, signal_928}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_931 ( .s (signal_745), .b ({signal_2582, signal_1847}), .a ({signal_2653, signal_1783}), .c ({signal_2924, signal_929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_934 ( .s (signal_404), .b ({signal_2560, signal_1838}), .a ({signal_2925, signal_932}), .c ({signal_3109, signal_931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_935 ( .s (signal_745), .b ({signal_2585, signal_1846}), .a ({signal_2656, signal_1782}), .c ({signal_2925, signal_932}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_938 ( .s (signal_404), .b ({signal_2563, signal_1509}), .a ({signal_2926, signal_935}), .c ({signal_3110, signal_934}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_939 ( .s (signal_745), .b ({signal_2588, signal_1837}), .a ({signal_2659, signal_1773}), .c ({signal_2926, signal_935}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_942 ( .s (signal_404), .b ({signal_2566, signal_1508}), .a ({signal_2927, signal_938}), .c ({signal_3111, signal_937}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_943 ( .s (signal_745), .b ({signal_2591, signal_1836}), .a ({signal_2662, signal_1772}), .c ({signal_2927, signal_938}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_946 ( .s (signal_404), .b ({signal_2569, signal_1507}), .a ({signal_2928, signal_941}), .c ({signal_3112, signal_940}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_947 ( .s (signal_745), .b ({signal_2594, signal_1835}), .a ({signal_2665, signal_1771}), .c ({signal_2928, signal_941}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_950 ( .s (signal_404), .b ({signal_2572, signal_1506}), .a ({signal_2929, signal_944}), .c ({signal_3113, signal_943}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_951 ( .s (signal_745), .b ({signal_2597, signal_1834}), .a ({signal_2668, signal_1770}), .c ({signal_2929, signal_944}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_954 ( .s (signal_404), .b ({signal_2575, signal_1505}), .a ({signal_2930, signal_947}), .c ({signal_3114, signal_946}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_955 ( .s (signal_745), .b ({signal_2600, signal_1833}), .a ({signal_2671, signal_1769}), .c ({signal_2930, signal_947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_958 ( .s (signal_404), .b ({signal_2578, signal_1504}), .a ({signal_2931, signal_950}), .c ({signal_3115, signal_949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_959 ( .s (signal_745), .b ({signal_2603, signal_1832}), .a ({signal_2674, signal_1768}), .c ({signal_2931, signal_950}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_962 ( .s (signal_404), .b ({signal_2581, signal_1503}), .a ({signal_2932, signal_953}), .c ({signal_3116, signal_952}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_963 ( .s (signal_745), .b ({signal_2606, signal_1831}), .a ({signal_2677, signal_1767}), .c ({signal_2932, signal_953}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_966 ( .s (signal_404), .b ({signal_2584, signal_1502}), .a ({signal_2933, signal_956}), .c ({signal_3117, signal_955}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_967 ( .s (signal_745), .b ({signal_2609, signal_1830}), .a ({signal_2680, signal_1766}), .c ({signal_2933, signal_956}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_970 ( .s (signal_754), .b ({signal_2587, signal_1821}), .a ({signal_2934, signal_959}), .c ({signal_3342, signal_958}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_971 ( .s (signal_746), .b ({signal_2612, signal_1829}), .a ({signal_2683, signal_1749}), .c ({signal_2934, signal_959}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_974 ( .s (signal_754), .b ({signal_2590, signal_1820}), .a ({signal_2935, signal_962}), .c ({signal_3343, signal_961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_975 ( .s (signal_746), .b ({signal_2615, signal_1828}), .a ({signal_2686, signal_1748}), .c ({signal_2935, signal_962}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_978 ( .s (signal_754), .b ({signal_2593, signal_1819}), .a ({signal_2936, signal_965}), .c ({signal_3344, signal_964}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_979 ( .s (signal_746), .b ({signal_2618, signal_1827}), .a ({signal_2689, signal_1747}), .c ({signal_2936, signal_965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_982 ( .s (signal_754), .b ({signal_2596, signal_1818}), .a ({signal_2937, signal_968}), .c ({signal_3345, signal_967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_983 ( .s (signal_746), .b ({signal_2621, signal_1826}), .a ({signal_2692, signal_1746}), .c ({signal_2937, signal_968}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_986 ( .s (signal_754), .b ({signal_2599, signal_1817}), .a ({signal_2938, signal_971}), .c ({signal_3346, signal_970}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_987 ( .s (signal_746), .b ({signal_2624, signal_1825}), .a ({signal_2695, signal_1745}), .c ({signal_2938, signal_971}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_990 ( .s (signal_754), .b ({signal_2602, signal_1816}), .a ({signal_2939, signal_974}), .c ({signal_3347, signal_973}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_991 ( .s (signal_746), .b ({signal_2627, signal_1824}), .a ({signal_2698, signal_1744}), .c ({signal_2939, signal_974}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_994 ( .s (signal_754), .b ({signal_2605, signal_1815}), .a ({signal_2940, signal_977}), .c ({signal_3348, signal_976}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_995 ( .s (signal_746), .b ({signal_2630, signal_1823}), .a ({signal_2701, signal_1743}), .c ({signal_2940, signal_977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_998 ( .s (signal_754), .b ({signal_2608, signal_1814}), .a ({signal_2941, signal_980}), .c ({signal_3349, signal_979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_999 ( .s (signal_746), .b ({signal_2633, signal_1822}), .a ({signal_2704, signal_1742}), .c ({signal_2941, signal_980}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1002 ( .s (signal_754), .b ({signal_2611, signal_1805}), .a ({signal_2942, signal_983}), .c ({signal_3350, signal_982}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1003 ( .s (signal_746), .b ({signal_2636, signal_1813}), .a ({signal_2707, signal_1733}), .c ({signal_2942, signal_983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1006 ( .s (signal_754), .b ({signal_2614, signal_1804}), .a ({signal_2943, signal_986}), .c ({signal_3351, signal_985}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1007 ( .s (signal_746), .b ({signal_2639, signal_1812}), .a ({signal_2710, signal_1732}), .c ({signal_2943, signal_986}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1010 ( .s (signal_754), .b ({signal_2617, signal_1803}), .a ({signal_2944, signal_989}), .c ({signal_3352, signal_988}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1011 ( .s (signal_746), .b ({signal_2642, signal_1811}), .a ({signal_2713, signal_1731}), .c ({signal_2944, signal_989}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1014 ( .s (signal_754), .b ({signal_2620, signal_1802}), .a ({signal_2945, signal_992}), .c ({signal_3353, signal_991}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1015 ( .s (signal_746), .b ({signal_2645, signal_1810}), .a ({signal_2716, signal_1730}), .c ({signal_2945, signal_992}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1018 ( .s (signal_754), .b ({signal_2623, signal_1801}), .a ({signal_2946, signal_995}), .c ({signal_3354, signal_994}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1019 ( .s (signal_746), .b ({signal_2648, signal_1809}), .a ({signal_2719, signal_1729}), .c ({signal_2946, signal_995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1022 ( .s (signal_754), .b ({signal_2626, signal_1800}), .a ({signal_2947, signal_998}), .c ({signal_3355, signal_997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1023 ( .s (signal_746), .b ({signal_2651, signal_1808}), .a ({signal_2722, signal_1728}), .c ({signal_2947, signal_998}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1026 ( .s (signal_754), .b ({signal_2629, signal_1799}), .a ({signal_2948, signal_1001}), .c ({signal_3356, signal_1000}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1027 ( .s (signal_746), .b ({signal_2654, signal_1807}), .a ({signal_2725, signal_1727}), .c ({signal_2948, signal_1001}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1030 ( .s (signal_754), .b ({signal_2632, signal_1798}), .a ({signal_2949, signal_1004}), .c ({signal_3357, signal_1003}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1031 ( .s (signal_746), .b ({signal_2657, signal_1806}), .a ({signal_2728, signal_1726}), .c ({signal_2949, signal_1004}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1034 ( .s (signal_755), .b ({signal_2635, signal_1789}), .a ({signal_2950, signal_1007}), .c ({signal_3358, signal_1006}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1035 ( .s (signal_747), .b ({signal_2660, signal_1797}), .a ({signal_2731, signal_1717}), .c ({signal_2950, signal_1007}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1038 ( .s (signal_755), .b ({signal_2638, signal_1788}), .a ({signal_2951, signal_1010}), .c ({signal_3359, signal_1009}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1039 ( .s (signal_747), .b ({signal_2663, signal_1796}), .a ({signal_2734, signal_1716}), .c ({signal_2951, signal_1010}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1042 ( .s (signal_755), .b ({signal_2641, signal_1787}), .a ({signal_2952, signal_1013}), .c ({signal_3360, signal_1012}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1043 ( .s (signal_747), .b ({signal_2666, signal_1795}), .a ({signal_2737, signal_1715}), .c ({signal_2952, signal_1013}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1046 ( .s (signal_755), .b ({signal_2644, signal_1786}), .a ({signal_2953, signal_1016}), .c ({signal_3361, signal_1015}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1047 ( .s (signal_747), .b ({signal_2669, signal_1794}), .a ({signal_2740, signal_1714}), .c ({signal_2953, signal_1016}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1050 ( .s (signal_755), .b ({signal_2647, signal_1785}), .a ({signal_2954, signal_1019}), .c ({signal_3362, signal_1018}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1051 ( .s (signal_747), .b ({signal_2672, signal_1793}), .a ({signal_2743, signal_1713}), .c ({signal_2954, signal_1019}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1054 ( .s (signal_755), .b ({signal_2650, signal_1784}), .a ({signal_2955, signal_1022}), .c ({signal_3363, signal_1021}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1055 ( .s (signal_747), .b ({signal_2675, signal_1792}), .a ({signal_2746, signal_1712}), .c ({signal_2955, signal_1022}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1058 ( .s (signal_755), .b ({signal_2653, signal_1783}), .a ({signal_2956, signal_1025}), .c ({signal_3364, signal_1024}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1059 ( .s (signal_747), .b ({signal_2678, signal_1791}), .a ({signal_2749, signal_1711}), .c ({signal_2956, signal_1025}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1062 ( .s (signal_755), .b ({signal_2656, signal_1782}), .a ({signal_2957, signal_1028}), .c ({signal_3365, signal_1027}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1063 ( .s (signal_747), .b ({signal_2681, signal_1790}), .a ({signal_2752, signal_1710}), .c ({signal_2957, signal_1028}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1066 ( .s (signal_755), .b ({signal_2659, signal_1773}), .a ({signal_2958, signal_1031}), .c ({signal_3366, signal_1030}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1067 ( .s (signal_747), .b ({signal_2684, signal_1781}), .a ({signal_2755, signal_1701}), .c ({signal_2958, signal_1031}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1070 ( .s (signal_755), .b ({signal_2662, signal_1772}), .a ({signal_2959, signal_1034}), .c ({signal_3367, signal_1033}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1071 ( .s (signal_747), .b ({signal_2687, signal_1780}), .a ({signal_2758, signal_1700}), .c ({signal_2959, signal_1034}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1074 ( .s (signal_755), .b ({signal_2665, signal_1771}), .a ({signal_2960, signal_1037}), .c ({signal_3368, signal_1036}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1075 ( .s (signal_747), .b ({signal_2690, signal_1779}), .a ({signal_2761, signal_1699}), .c ({signal_2960, signal_1037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1078 ( .s (signal_755), .b ({signal_2668, signal_1770}), .a ({signal_2961, signal_1040}), .c ({signal_3369, signal_1039}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1079 ( .s (signal_747), .b ({signal_2693, signal_1778}), .a ({signal_2764, signal_1698}), .c ({signal_2961, signal_1040}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1082 ( .s (signal_755), .b ({signal_2671, signal_1769}), .a ({signal_2962, signal_1043}), .c ({signal_3370, signal_1042}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1083 ( .s (signal_747), .b ({signal_2696, signal_1777}), .a ({signal_2767, signal_1697}), .c ({signal_2962, signal_1043}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1086 ( .s (signal_755), .b ({signal_2674, signal_1768}), .a ({signal_2963, signal_1046}), .c ({signal_3371, signal_1045}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1087 ( .s (signal_747), .b ({signal_2699, signal_1776}), .a ({signal_2770, signal_1696}), .c ({signal_2963, signal_1046}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1090 ( .s (signal_755), .b ({signal_2677, signal_1767}), .a ({signal_2964, signal_1049}), .c ({signal_3372, signal_1048}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1091 ( .s (signal_747), .b ({signal_2702, signal_1775}), .a ({signal_2773, signal_1695}), .c ({signal_2964, signal_1049}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1094 ( .s (signal_755), .b ({signal_2680, signal_1766}), .a ({signal_2965, signal_1052}), .c ({signal_3373, signal_1051}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1095 ( .s (signal_747), .b ({signal_2705, signal_1774}), .a ({signal_2776, signal_1694}), .c ({signal_2965, signal_1052}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1130 ( .s (signal_756), .b ({signal_2707, signal_1733}), .a ({signal_2966, signal_1079}), .c ({signal_3382, signal_1078}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1131 ( .s (signal_748), .b ({signal_2732, signal_1741}), .a ({signal_2020, signal_758}), .c ({signal_2966, signal_1079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1134 ( .s (signal_756), .b ({signal_2710, signal_1732}), .a ({signal_2967, signal_1082}), .c ({signal_3383, signal_1081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1135 ( .s (signal_748), .b ({signal_2735, signal_1740}), .a ({signal_2018, signal_759}), .c ({signal_2967, signal_1082}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1138 ( .s (signal_756), .b ({signal_2713, signal_1731}), .a ({signal_2968, signal_1085}), .c ({signal_3384, signal_1084}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1139 ( .s (signal_748), .b ({signal_2738, signal_1739}), .a ({signal_2016, signal_760}), .c ({signal_2968, signal_1085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1142 ( .s (signal_756), .b ({signal_2716, signal_1730}), .a ({signal_2969, signal_1088}), .c ({signal_3385, signal_1087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1143 ( .s (signal_748), .b ({signal_2741, signal_1738}), .a ({signal_2014, signal_761}), .c ({signal_2969, signal_1088}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1146 ( .s (signal_756), .b ({signal_2719, signal_1729}), .a ({signal_2970, signal_1091}), .c ({signal_3386, signal_1090}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1147 ( .s (signal_748), .b ({signal_2744, signal_1737}), .a ({signal_2012, signal_762}), .c ({signal_2970, signal_1091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1150 ( .s (signal_756), .b ({signal_2722, signal_1728}), .a ({signal_2971, signal_1094}), .c ({signal_3387, signal_1093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1151 ( .s (signal_748), .b ({signal_2747, signal_1736}), .a ({signal_2010, signal_763}), .c ({signal_2971, signal_1094}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1154 ( .s (signal_756), .b ({signal_2725, signal_1727}), .a ({signal_2972, signal_1097}), .c ({signal_3388, signal_1096}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1155 ( .s (signal_748), .b ({signal_2750, signal_1735}), .a ({signal_2008, signal_764}), .c ({signal_2972, signal_1097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1158 ( .s (signal_756), .b ({signal_2728, signal_1726}), .a ({signal_2973, signal_1100}), .c ({signal_3389, signal_1099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1159 ( .s (signal_748), .b ({signal_2753, signal_1734}), .a ({signal_2006, signal_765}), .c ({signal_2973, signal_1100}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1162 ( .s (signal_757), .b ({signal_2731, signal_1717}), .a ({signal_2974, signal_1103}), .c ({signal_3390, signal_1102}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1163 ( .s (signal_749), .b ({signal_2756, signal_1725}), .a ({signal_2443, signal_1909}), .c ({signal_2974, signal_1103}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1166 ( .s (signal_757), .b ({signal_2734, signal_1716}), .a ({signal_2975, signal_1106}), .c ({signal_3391, signal_1105}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1167 ( .s (signal_749), .b ({signal_2759, signal_1724}), .a ({signal_2446, signal_1908}), .c ({signal_2975, signal_1106}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1170 ( .s (signal_757), .b ({signal_2737, signal_1715}), .a ({signal_2976, signal_1109}), .c ({signal_3392, signal_1108}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1171 ( .s (signal_749), .b ({signal_2762, signal_1723}), .a ({signal_2449, signal_1907}), .c ({signal_2976, signal_1109}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1174 ( .s (signal_757), .b ({signal_2740, signal_1714}), .a ({signal_2977, signal_1112}), .c ({signal_3393, signal_1111}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1175 ( .s (signal_749), .b ({signal_2765, signal_1722}), .a ({signal_2452, signal_1906}), .c ({signal_2977, signal_1112}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1178 ( .s (signal_757), .b ({signal_2743, signal_1713}), .a ({signal_2978, signal_1115}), .c ({signal_3394, signal_1114}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1179 ( .s (signal_749), .b ({signal_2768, signal_1721}), .a ({signal_2455, signal_1905}), .c ({signal_2978, signal_1115}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1182 ( .s (signal_757), .b ({signal_2746, signal_1712}), .a ({signal_2979, signal_1118}), .c ({signal_3395, signal_1117}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1183 ( .s (signal_749), .b ({signal_2771, signal_1720}), .a ({signal_2458, signal_1904}), .c ({signal_2979, signal_1118}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1186 ( .s (signal_757), .b ({signal_2749, signal_1711}), .a ({signal_2980, signal_1121}), .c ({signal_3396, signal_1120}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1187 ( .s (signal_749), .b ({signal_2774, signal_1719}), .a ({signal_2461, signal_1903}), .c ({signal_2980, signal_1121}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1190 ( .s (signal_757), .b ({signal_2752, signal_1710}), .a ({signal_2981, signal_1124}), .c ({signal_3397, signal_1123}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1191 ( .s (signal_749), .b ({signal_2777, signal_1718}), .a ({signal_2464, signal_1902}), .c ({signal_2981, signal_1124}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1194 ( .s (signal_757), .b ({signal_2755, signal_1701}), .a ({signal_2982, signal_1127}), .c ({signal_3398, signal_1126}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1195 ( .s (signal_749), .b ({signal_2779, signal_1709}), .a ({signal_2467, signal_1893}), .c ({signal_2982, signal_1127}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1198 ( .s (signal_757), .b ({signal_2758, signal_1700}), .a ({signal_2983, signal_1130}), .c ({signal_3399, signal_1129}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1199 ( .s (signal_749), .b ({signal_2781, signal_1708}), .a ({signal_2470, signal_1892}), .c ({signal_2983, signal_1130}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1202 ( .s (signal_757), .b ({signal_2761, signal_1699}), .a ({signal_2984, signal_1133}), .c ({signal_3400, signal_1132}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1203 ( .s (signal_749), .b ({signal_2783, signal_1707}), .a ({signal_2473, signal_1891}), .c ({signal_2984, signal_1133}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1206 ( .s (signal_757), .b ({signal_2764, signal_1698}), .a ({signal_2985, signal_1136}), .c ({signal_3401, signal_1135}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1207 ( .s (signal_749), .b ({signal_2785, signal_1706}), .a ({signal_2476, signal_1890}), .c ({signal_2985, signal_1136}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1210 ( .s (signal_757), .b ({signal_2767, signal_1697}), .a ({signal_2986, signal_1139}), .c ({signal_3402, signal_1138}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1211 ( .s (signal_749), .b ({signal_2787, signal_1705}), .a ({signal_2479, signal_1889}), .c ({signal_2986, signal_1139}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1214 ( .s (signal_757), .b ({signal_2770, signal_1696}), .a ({signal_2987, signal_1142}), .c ({signal_3403, signal_1141}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1215 ( .s (signal_749), .b ({signal_2789, signal_1704}), .a ({signal_2482, signal_1888}), .c ({signal_2987, signal_1142}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1218 ( .s (signal_757), .b ({signal_2773, signal_1695}), .a ({signal_2988, signal_1145}), .c ({signal_3404, signal_1144}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1219 ( .s (signal_749), .b ({signal_2791, signal_1703}), .a ({signal_2485, signal_1887}), .c ({signal_2988, signal_1145}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1222 ( .s (signal_757), .b ({signal_2776, signal_1694}), .a ({signal_2989, signal_1148}), .c ({signal_3405, signal_1147}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1223 ( .s (signal_749), .b ({signal_2793, signal_1702}), .a ({signal_2488, signal_1886}), .c ({signal_2989, signal_1148}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1226 ( .s (signal_400), .b ({signal_2020, signal_758}), .a ({signal_2021, signal_1693}), .c ({signal_3118, signal_1685}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1227 ( .s (signal_400), .b ({signal_2018, signal_759}), .a ({signal_2019, signal_1692}), .c ({signal_3119, signal_1684}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1228 ( .s (signal_400), .b ({signal_2016, signal_760}), .a ({signal_2017, signal_1691}), .c ({signal_3120, signal_1683}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1229 ( .s (signal_400), .b ({signal_2014, signal_761}), .a ({signal_2015, signal_1690}), .c ({signal_3121, signal_1682}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1230 ( .s (signal_400), .b ({signal_2012, signal_762}), .a ({signal_2013, signal_1689}), .c ({signal_3122, signal_1681}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1231 ( .s (signal_400), .b ({signal_2010, signal_763}), .a ({signal_2011, signal_1688}), .c ({signal_3123, signal_1680}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1232 ( .s (signal_400), .b ({signal_2008, signal_764}), .a ({signal_2009, signal_1687}), .c ({signal_3124, signal_1679}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1233 ( .s (signal_400), .b ({signal_2006, signal_765}), .a ({signal_2007, signal_1686}), .c ({signal_3125, signal_1678}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1234 ( .s (signal_733), .b ({key_s1[120], key_s0[120]}), .a ({signal_3118, signal_1685}), .c ({signal_3271, signal_1933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1235 ( .s (signal_733), .b ({key_s1[121], key_s0[121]}), .a ({signal_3119, signal_1684}), .c ({signal_3273, signal_1932}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1236 ( .s (signal_733), .b ({key_s1[122], key_s0[122]}), .a ({signal_3120, signal_1683}), .c ({signal_3275, signal_1931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1237 ( .s (signal_733), .b ({key_s1[123], key_s0[123]}), .a ({signal_3121, signal_1682}), .c ({signal_3277, signal_1930}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1238 ( .s (signal_733), .b ({key_s1[124], key_s0[124]}), .a ({signal_3122, signal_1681}), .c ({signal_3279, signal_1929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1239 ( .s (signal_733), .b ({key_s1[125], key_s0[125]}), .a ({signal_3123, signal_1680}), .c ({signal_3281, signal_1928}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1240 ( .s (signal_733), .b ({key_s1[126], key_s0[126]}), .a ({signal_3124, signal_1679}), .c ({signal_3283, signal_1927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1241 ( .s (signal_733), .b ({key_s1[127], key_s0[127]}), .a ({signal_3125, signal_1678}), .c ({signal_3285, signal_1926}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1242 ( .s (signal_733), .b ({key_s1[112], key_s0[112]}), .a ({signal_2443, signal_1909}), .c ({signal_2444, signal_1925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1243 ( .s (signal_733), .b ({key_s1[113], key_s0[113]}), .a ({signal_2446, signal_1908}), .c ({signal_2447, signal_1924}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1244 ( .s (signal_733), .b ({key_s1[114], key_s0[114]}), .a ({signal_2449, signal_1907}), .c ({signal_2450, signal_1923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1245 ( .s (signal_733), .b ({key_s1[115], key_s0[115]}), .a ({signal_2452, signal_1906}), .c ({signal_2453, signal_1922}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1246 ( .s (signal_733), .b ({key_s1[116], key_s0[116]}), .a ({signal_2455, signal_1905}), .c ({signal_2456, signal_1921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1247 ( .s (signal_733), .b ({key_s1[117], key_s0[117]}), .a ({signal_2458, signal_1904}), .c ({signal_2459, signal_1920}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1248 ( .s (signal_733), .b ({key_s1[118], key_s0[118]}), .a ({signal_2461, signal_1903}), .c ({signal_2462, signal_1919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1249 ( .s (signal_733), .b ({key_s1[119], key_s0[119]}), .a ({signal_2464, signal_1902}), .c ({signal_2465, signal_1918}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1250 ( .s (signal_734), .b ({key_s1[104], key_s0[104]}), .a ({signal_2467, signal_1893}), .c ({signal_2468, signal_1917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1251 ( .s (signal_734), .b ({key_s1[105], key_s0[105]}), .a ({signal_2470, signal_1892}), .c ({signal_2471, signal_1916}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1252 ( .s (signal_734), .b ({key_s1[106], key_s0[106]}), .a ({signal_2473, signal_1891}), .c ({signal_2474, signal_1915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1253 ( .s (signal_734), .b ({key_s1[107], key_s0[107]}), .a ({signal_2476, signal_1890}), .c ({signal_2477, signal_1914}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1254 ( .s (signal_734), .b ({key_s1[108], key_s0[108]}), .a ({signal_2479, signal_1889}), .c ({signal_2480, signal_1913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1255 ( .s (signal_734), .b ({key_s1[109], key_s0[109]}), .a ({signal_2482, signal_1888}), .c ({signal_2483, signal_1912}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1256 ( .s (signal_734), .b ({key_s1[110], key_s0[110]}), .a ({signal_2485, signal_1887}), .c ({signal_2486, signal_1911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1257 ( .s (signal_734), .b ({key_s1[111], key_s0[111]}), .a ({signal_2488, signal_1886}), .c ({signal_2489, signal_1910}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1258 ( .s (signal_734), .b ({key_s1[96], key_s0[96]}), .a ({signal_2491, signal_1877}), .c ({signal_2492, signal_1901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1259 ( .s (signal_734), .b ({key_s1[97], key_s0[97]}), .a ({signal_2494, signal_1876}), .c ({signal_2495, signal_1900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1260 ( .s (signal_734), .b ({key_s1[98], key_s0[98]}), .a ({signal_2497, signal_1875}), .c ({signal_2498, signal_1899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1261 ( .s (signal_734), .b ({key_s1[99], key_s0[99]}), .a ({signal_2500, signal_1874}), .c ({signal_2501, signal_1898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1262 ( .s (signal_734), .b ({key_s1[100], key_s0[100]}), .a ({signal_2503, signal_1873}), .c ({signal_2504, signal_1897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1263 ( .s (signal_734), .b ({key_s1[101], key_s0[101]}), .a ({signal_2506, signal_1872}), .c ({signal_2507, signal_1896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1264 ( .s (signal_734), .b ({key_s1[102], key_s0[102]}), .a ({signal_2509, signal_1871}), .c ({signal_2510, signal_1895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1265 ( .s (signal_734), .b ({key_s1[103], key_s0[103]}), .a ({signal_2512, signal_1870}), .c ({signal_2513, signal_1894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1266 ( .s (signal_735), .b ({key_s1[88], key_s0[88]}), .a ({signal_2515, signal_1861}), .c ({signal_2516, signal_1885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1267 ( .s (signal_735), .b ({key_s1[89], key_s0[89]}), .a ({signal_2518, signal_1860}), .c ({signal_2519, signal_1884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1268 ( .s (signal_735), .b ({key_s1[90], key_s0[90]}), .a ({signal_2521, signal_1859}), .c ({signal_2522, signal_1883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1269 ( .s (signal_735), .b ({key_s1[91], key_s0[91]}), .a ({signal_2524, signal_1858}), .c ({signal_2525, signal_1882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1270 ( .s (signal_735), .b ({key_s1[92], key_s0[92]}), .a ({signal_2527, signal_1857}), .c ({signal_2528, signal_1881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1271 ( .s (signal_735), .b ({key_s1[93], key_s0[93]}), .a ({signal_2530, signal_1856}), .c ({signal_2531, signal_1880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1272 ( .s (signal_735), .b ({key_s1[94], key_s0[94]}), .a ({signal_2533, signal_1855}), .c ({signal_2534, signal_1879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1273 ( .s (signal_735), .b ({key_s1[95], key_s0[95]}), .a ({signal_2536, signal_1854}), .c ({signal_2537, signal_1878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1274 ( .s (signal_735), .b ({key_s1[80], key_s0[80]}), .a ({signal_2539, signal_1845}), .c ({signal_2540, signal_1869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1275 ( .s (signal_735), .b ({key_s1[81], key_s0[81]}), .a ({signal_2542, signal_1844}), .c ({signal_2543, signal_1868}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1276 ( .s (signal_735), .b ({key_s1[82], key_s0[82]}), .a ({signal_2545, signal_1843}), .c ({signal_2546, signal_1867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1277 ( .s (signal_735), .b ({key_s1[83], key_s0[83]}), .a ({signal_2548, signal_1842}), .c ({signal_2549, signal_1866}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1278 ( .s (signal_735), .b ({key_s1[84], key_s0[84]}), .a ({signal_2551, signal_1841}), .c ({signal_2552, signal_1865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1279 ( .s (signal_735), .b ({key_s1[85], key_s0[85]}), .a ({signal_2554, signal_1840}), .c ({signal_2555, signal_1864}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1280 ( .s (signal_735), .b ({key_s1[86], key_s0[86]}), .a ({signal_2557, signal_1839}), .c ({signal_2558, signal_1863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1281 ( .s (signal_735), .b ({key_s1[87], key_s0[87]}), .a ({signal_2560, signal_1838}), .c ({signal_2561, signal_1862}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1282 ( .s (signal_736), .b ({key_s1[72], key_s0[72]}), .a ({signal_2563, signal_1509}), .c ({signal_2564, signal_1853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1283 ( .s (signal_736), .b ({key_s1[73], key_s0[73]}), .a ({signal_2566, signal_1508}), .c ({signal_2567, signal_1852}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1284 ( .s (signal_736), .b ({key_s1[74], key_s0[74]}), .a ({signal_2569, signal_1507}), .c ({signal_2570, signal_1851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1285 ( .s (signal_736), .b ({key_s1[75], key_s0[75]}), .a ({signal_2572, signal_1506}), .c ({signal_2573, signal_1850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1286 ( .s (signal_736), .b ({key_s1[76], key_s0[76]}), .a ({signal_2575, signal_1505}), .c ({signal_2576, signal_1849}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1287 ( .s (signal_736), .b ({key_s1[77], key_s0[77]}), .a ({signal_2578, signal_1504}), .c ({signal_2579, signal_1848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1288 ( .s (signal_736), .b ({key_s1[78], key_s0[78]}), .a ({signal_2581, signal_1503}), .c ({signal_2582, signal_1847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1289 ( .s (signal_736), .b ({key_s1[79], key_s0[79]}), .a ({signal_2584, signal_1502}), .c ({signal_2585, signal_1846}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1290 ( .s (signal_736), .b ({key_s1[64], key_s0[64]}), .a ({signal_2587, signal_1821}), .c ({signal_2588, signal_1837}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1291 ( .s (signal_736), .b ({key_s1[65], key_s0[65]}), .a ({signal_2590, signal_1820}), .c ({signal_2591, signal_1836}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1292 ( .s (signal_736), .b ({key_s1[66], key_s0[66]}), .a ({signal_2593, signal_1819}), .c ({signal_2594, signal_1835}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1293 ( .s (signal_736), .b ({key_s1[67], key_s0[67]}), .a ({signal_2596, signal_1818}), .c ({signal_2597, signal_1834}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1294 ( .s (signal_736), .b ({key_s1[68], key_s0[68]}), .a ({signal_2599, signal_1817}), .c ({signal_2600, signal_1833}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1295 ( .s (signal_736), .b ({key_s1[69], key_s0[69]}), .a ({signal_2602, signal_1816}), .c ({signal_2603, signal_1832}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1296 ( .s (signal_736), .b ({key_s1[70], key_s0[70]}), .a ({signal_2605, signal_1815}), .c ({signal_2606, signal_1831}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1297 ( .s (signal_736), .b ({key_s1[71], key_s0[71]}), .a ({signal_2608, signal_1814}), .c ({signal_2609, signal_1830}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1298 ( .s (signal_737), .b ({key_s1[56], key_s0[56]}), .a ({signal_2611, signal_1805}), .c ({signal_2612, signal_1829}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1299 ( .s (signal_737), .b ({key_s1[57], key_s0[57]}), .a ({signal_2614, signal_1804}), .c ({signal_2615, signal_1828}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1300 ( .s (signal_737), .b ({key_s1[58], key_s0[58]}), .a ({signal_2617, signal_1803}), .c ({signal_2618, signal_1827}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1301 ( .s (signal_737), .b ({key_s1[59], key_s0[59]}), .a ({signal_2620, signal_1802}), .c ({signal_2621, signal_1826}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1302 ( .s (signal_737), .b ({key_s1[60], key_s0[60]}), .a ({signal_2623, signal_1801}), .c ({signal_2624, signal_1825}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1303 ( .s (signal_737), .b ({key_s1[61], key_s0[61]}), .a ({signal_2626, signal_1800}), .c ({signal_2627, signal_1824}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1304 ( .s (signal_737), .b ({key_s1[62], key_s0[62]}), .a ({signal_2629, signal_1799}), .c ({signal_2630, signal_1823}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1305 ( .s (signal_737), .b ({key_s1[63], key_s0[63]}), .a ({signal_2632, signal_1798}), .c ({signal_2633, signal_1822}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1306 ( .s (signal_737), .b ({key_s1[48], key_s0[48]}), .a ({signal_2635, signal_1789}), .c ({signal_2636, signal_1813}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1307 ( .s (signal_737), .b ({key_s1[49], key_s0[49]}), .a ({signal_2638, signal_1788}), .c ({signal_2639, signal_1812}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1308 ( .s (signal_737), .b ({key_s1[50], key_s0[50]}), .a ({signal_2641, signal_1787}), .c ({signal_2642, signal_1811}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1309 ( .s (signal_737), .b ({key_s1[51], key_s0[51]}), .a ({signal_2644, signal_1786}), .c ({signal_2645, signal_1810}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1310 ( .s (signal_737), .b ({key_s1[52], key_s0[52]}), .a ({signal_2647, signal_1785}), .c ({signal_2648, signal_1809}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1311 ( .s (signal_737), .b ({key_s1[53], key_s0[53]}), .a ({signal_2650, signal_1784}), .c ({signal_2651, signal_1808}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1312 ( .s (signal_737), .b ({key_s1[54], key_s0[54]}), .a ({signal_2653, signal_1783}), .c ({signal_2654, signal_1807}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1313 ( .s (signal_737), .b ({key_s1[55], key_s0[55]}), .a ({signal_2656, signal_1782}), .c ({signal_2657, signal_1806}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1314 ( .s (signal_738), .b ({key_s1[40], key_s0[40]}), .a ({signal_2659, signal_1773}), .c ({signal_2660, signal_1797}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1315 ( .s (signal_738), .b ({key_s1[41], key_s0[41]}), .a ({signal_2662, signal_1772}), .c ({signal_2663, signal_1796}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1316 ( .s (signal_738), .b ({key_s1[42], key_s0[42]}), .a ({signal_2665, signal_1771}), .c ({signal_2666, signal_1795}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1317 ( .s (signal_738), .b ({key_s1[43], key_s0[43]}), .a ({signal_2668, signal_1770}), .c ({signal_2669, signal_1794}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1318 ( .s (signal_738), .b ({key_s1[44], key_s0[44]}), .a ({signal_2671, signal_1769}), .c ({signal_2672, signal_1793}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1319 ( .s (signal_738), .b ({key_s1[45], key_s0[45]}), .a ({signal_2674, signal_1768}), .c ({signal_2675, signal_1792}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1320 ( .s (signal_738), .b ({key_s1[46], key_s0[46]}), .a ({signal_2677, signal_1767}), .c ({signal_2678, signal_1791}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1321 ( .s (signal_738), .b ({key_s1[47], key_s0[47]}), .a ({signal_2680, signal_1766}), .c ({signal_2681, signal_1790}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1322 ( .s (signal_738), .b ({key_s1[32], key_s0[32]}), .a ({signal_2683, signal_1749}), .c ({signal_2684, signal_1781}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1323 ( .s (signal_738), .b ({key_s1[33], key_s0[33]}), .a ({signal_2686, signal_1748}), .c ({signal_2687, signal_1780}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1324 ( .s (signal_738), .b ({key_s1[34], key_s0[34]}), .a ({signal_2689, signal_1747}), .c ({signal_2690, signal_1779}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1325 ( .s (signal_738), .b ({key_s1[35], key_s0[35]}), .a ({signal_2692, signal_1746}), .c ({signal_2693, signal_1778}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1326 ( .s (signal_738), .b ({key_s1[36], key_s0[36]}), .a ({signal_2695, signal_1745}), .c ({signal_2696, signal_1777}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1327 ( .s (signal_738), .b ({key_s1[37], key_s0[37]}), .a ({signal_2698, signal_1744}), .c ({signal_2699, signal_1776}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1328 ( .s (signal_738), .b ({key_s1[38], key_s0[38]}), .a ({signal_2701, signal_1743}), .c ({signal_2702, signal_1775}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1329 ( .s (signal_738), .b ({key_s1[39], key_s0[39]}), .a ({signal_2704, signal_1742}), .c ({signal_2705, signal_1774}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1330 ( .s (signal_739), .b ({key_s1[24], key_s0[24]}), .a ({signal_2707, signal_1733}), .c ({signal_2708, signal_1765}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1331 ( .s (signal_739), .b ({key_s1[25], key_s0[25]}), .a ({signal_2710, signal_1732}), .c ({signal_2711, signal_1764}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1332 ( .s (signal_739), .b ({key_s1[26], key_s0[26]}), .a ({signal_2713, signal_1731}), .c ({signal_2714, signal_1763}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1333 ( .s (signal_739), .b ({key_s1[27], key_s0[27]}), .a ({signal_2716, signal_1730}), .c ({signal_2717, signal_1762}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1334 ( .s (signal_739), .b ({key_s1[28], key_s0[28]}), .a ({signal_2719, signal_1729}), .c ({signal_2720, signal_1761}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1335 ( .s (signal_739), .b ({key_s1[29], key_s0[29]}), .a ({signal_2722, signal_1728}), .c ({signal_2723, signal_1760}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1336 ( .s (signal_739), .b ({key_s1[30], key_s0[30]}), .a ({signal_2725, signal_1727}), .c ({signal_2726, signal_1759}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1337 ( .s (signal_739), .b ({key_s1[31], key_s0[31]}), .a ({signal_2728, signal_1726}), .c ({signal_2729, signal_1758}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1338 ( .s (signal_739), .b ({key_s1[16], key_s0[16]}), .a ({signal_2731, signal_1717}), .c ({signal_2732, signal_1741}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1339 ( .s (signal_739), .b ({key_s1[17], key_s0[17]}), .a ({signal_2734, signal_1716}), .c ({signal_2735, signal_1740}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1340 ( .s (signal_739), .b ({key_s1[18], key_s0[18]}), .a ({signal_2737, signal_1715}), .c ({signal_2738, signal_1739}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1341 ( .s (signal_739), .b ({key_s1[19], key_s0[19]}), .a ({signal_2740, signal_1714}), .c ({signal_2741, signal_1738}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1342 ( .s (signal_739), .b ({key_s1[20], key_s0[20]}), .a ({signal_2743, signal_1713}), .c ({signal_2744, signal_1737}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1343 ( .s (signal_739), .b ({key_s1[21], key_s0[21]}), .a ({signal_2746, signal_1712}), .c ({signal_2747, signal_1736}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1344 ( .s (signal_739), .b ({key_s1[22], key_s0[22]}), .a ({signal_2749, signal_1711}), .c ({signal_2750, signal_1735}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1345 ( .s (signal_739), .b ({key_s1[23], key_s0[23]}), .a ({signal_2752, signal_1710}), .c ({signal_2753, signal_1734}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1346 ( .s (signal_740), .b ({key_s1[8], key_s0[8]}), .a ({signal_2755, signal_1701}), .c ({signal_2756, signal_1725}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1347 ( .s (signal_740), .b ({key_s1[9], key_s0[9]}), .a ({signal_2758, signal_1700}), .c ({signal_2759, signal_1724}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1348 ( .s (signal_740), .b ({key_s1[10], key_s0[10]}), .a ({signal_2761, signal_1699}), .c ({signal_2762, signal_1723}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1349 ( .s (signal_740), .b ({key_s1[11], key_s0[11]}), .a ({signal_2764, signal_1698}), .c ({signal_2765, signal_1722}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1350 ( .s (signal_740), .b ({key_s1[12], key_s0[12]}), .a ({signal_2767, signal_1697}), .c ({signal_2768, signal_1721}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1351 ( .s (signal_740), .b ({key_s1[13], key_s0[13]}), .a ({signal_2770, signal_1696}), .c ({signal_2771, signal_1720}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1352 ( .s (signal_740), .b ({key_s1[14], key_s0[14]}), .a ({signal_2773, signal_1695}), .c ({signal_2774, signal_1719}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1353 ( .s (signal_740), .b ({key_s1[15], key_s0[15]}), .a ({signal_2776, signal_1694}), .c ({signal_2777, signal_1718}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1354 ( .s (signal_740), .b ({key_s1[0], key_s0[0]}), .a ({signal_1983, signal_1493}), .c ({signal_2779, signal_1709}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1355 ( .s (signal_740), .b ({key_s1[1], key_s0[1]}), .a ({signal_1986, signal_1492}), .c ({signal_2781, signal_1708}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1356 ( .s (signal_740), .b ({key_s1[2], key_s0[2]}), .a ({signal_1989, signal_1491}), .c ({signal_2783, signal_1707}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1357 ( .s (signal_740), .b ({key_s1[3], key_s0[3]}), .a ({signal_1992, signal_1490}), .c ({signal_2785, signal_1706}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1358 ( .s (signal_740), .b ({key_s1[4], key_s0[4]}), .a ({signal_1995, signal_1489}), .c ({signal_2787, signal_1705}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1359 ( .s (signal_740), .b ({key_s1[5], key_s0[5]}), .a ({signal_1998, signal_1488}), .c ({signal_2789, signal_1704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1360 ( .s (signal_740), .b ({key_s1[6], key_s0[6]}), .a ({signal_2001, signal_1487}), .c ({signal_2791, signal_1703}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1361 ( .s (signal_740), .b ({key_s1[7], key_s0[7]}), .a ({signal_2004, signal_1486}), .c ({signal_2793, signal_1702}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1362 ( .a ({signal_2122, signal_1150}), .b ({signal_2024, signal_1151}), .c ({signal_2794, signal_1454}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1363 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2024, signal_1151}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1364 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2051, signal_1934}), .c ({signal_2122, signal_1150}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1365 ( .a ({signal_2123, signal_1152}), .b ({signal_2027, signal_1153}), .c ({signal_2795, signal_1455}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1366 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2027, signal_1153}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1367 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2053, signal_1935}), .c ({signal_2123, signal_1152}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1368 ( .a ({signal_2124, signal_1154}), .b ({signal_2030, signal_1155}), .c ({signal_2796, signal_1456}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1369 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2030, signal_1155}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1370 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2055, signal_1936}), .c ({signal_2124, signal_1154}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1371 ( .a ({signal_2797, signal_1156}), .b ({signal_2033, signal_1157}), .c ({signal_2838, signal_1457}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1372 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2033, signal_1157}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1373 ( .a ({signal_2046, signal_1942}), .b ({signal_2127, signal_1937}), .c ({signal_2797, signal_1156}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1374 ( .a ({signal_2798, signal_1158}), .b ({signal_2036, signal_1159}), .c ({signal_2839, signal_1458}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1375 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2036, signal_1159}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1376 ( .a ({signal_2047, signal_1943}), .b ({signal_2128, signal_1938}), .c ({signal_2798, signal_1158}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1377 ( .a ({signal_2125, signal_1160}), .b ({signal_2039, signal_1161}), .c ({signal_2799, signal_1459}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1378 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2039, signal_1161}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1379 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2058, signal_1939}), .c ({signal_2125, signal_1160}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1380 ( .a ({signal_2800, signal_1162}), .b ({signal_2042, signal_1163}), .c ({signal_2840, signal_1460}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1381 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2042, signal_1163}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1382 ( .a ({signal_2048, signal_1945}), .b ({signal_2129, signal_1940}), .c ({signal_2800, signal_1162}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1383 ( .a ({signal_2126, signal_1164}), .b ({signal_2045, signal_1165}), .c ({signal_2801, signal_1461}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1384 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2045, signal_1165}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1385 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2060, signal_1941}), .c ({signal_2126, signal_1164}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1386 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2046, signal_1942}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1387 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2047, signal_1943}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1388 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2048, signal_1945}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1389 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2051, signal_1934}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1390 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2053, signal_1935}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1391 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2055, signal_1936}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1392 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2062, signal_1946}), .c ({signal_2127, signal_1937}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1393 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2063, signal_1947}), .c ({signal_2128, signal_1938}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1394 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2058, signal_1939}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1395 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2064, signal_1949}), .c ({signal_2129, signal_1940}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1396 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2060, signal_1941}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1397 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2062, signal_1946}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1398 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2063, signal_1947}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1399 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2064, signal_1949}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1400 ( .a ({signal_2130, signal_1166}), .b ({signal_2065, signal_1167}), .c ({signal_2802, signal_1462}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1401 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2065, signal_1167}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1402 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2076, signal_1950}), .c ({signal_2130, signal_1166}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1403 ( .a ({signal_2131, signal_1168}), .b ({signal_2066, signal_1169}), .c ({signal_2803, signal_1463}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1404 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2066, signal_1169}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1405 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2077, signal_1951}), .c ({signal_2131, signal_1168}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1406 ( .a ({signal_2132, signal_1170}), .b ({signal_2067, signal_1171}), .c ({signal_2804, signal_1464}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1407 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2067, signal_1171}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1408 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2078, signal_1952}), .c ({signal_2132, signal_1170}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1409 ( .a ({signal_2805, signal_1172}), .b ({signal_2068, signal_1173}), .c ({signal_2841, signal_1465}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1410 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2068, signal_1173}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1411 ( .a ({signal_2073, signal_1184}), .b ({signal_2135, signal_1953}), .c ({signal_2805, signal_1172}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1412 ( .a ({signal_2806, signal_1174}), .b ({signal_2069, signal_1175}), .c ({signal_2842, signal_1466}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1413 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2069, signal_1175}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1414 ( .a ({signal_2074, signal_1183}), .b ({signal_2136, signal_1954}), .c ({signal_2806, signal_1174}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1415 ( .a ({signal_2133, signal_1176}), .b ({signal_2070, signal_1177}), .c ({signal_2807, signal_1467}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1416 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2070, signal_1177}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1417 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2079, signal_1955}), .c ({signal_2133, signal_1176}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1418 ( .a ({signal_2808, signal_1178}), .b ({signal_2071, signal_1179}), .c ({signal_2843, signal_1468}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1419 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2071, signal_1179}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1420 ( .a ({signal_2075, signal_1182}), .b ({signal_2137, signal_1956}), .c ({signal_2808, signal_1178}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1421 ( .a ({signal_2134, signal_1180}), .b ({signal_2072, signal_1181}), .c ({signal_2809, signal_1469}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1422 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2072, signal_1181}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1423 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2080, signal_1957}), .c ({signal_2134, signal_1180}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1424 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2073, signal_1184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1425 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2074, signal_1183}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1426 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2075, signal_1182}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1427 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2076, signal_1950}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1428 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2077, signal_1951}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1429 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2078, signal_1952}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1430 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2081, signal_1958}), .c ({signal_2135, signal_1953}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1431 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2082, signal_1959}), .c ({signal_2136, signal_1954}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1432 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2079, signal_1955}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1433 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2083, signal_1961}), .c ({signal_2137, signal_1956}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1434 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2080, signal_1957}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1435 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2081, signal_1958}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1436 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2082, signal_1959}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1437 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2083, signal_1961}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1438 ( .a ({signal_2138, signal_1185}), .b ({signal_2084, signal_1186}), .c ({signal_2810, signal_1470}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1439 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2084, signal_1186}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1440 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2095, signal_1962}), .c ({signal_2138, signal_1185}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1441 ( .a ({signal_2139, signal_1187}), .b ({signal_2085, signal_1188}), .c ({signal_2811, signal_1471}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1442 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2085, signal_1188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1443 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2096, signal_1963}), .c ({signal_2139, signal_1187}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1444 ( .a ({signal_2140, signal_1189}), .b ({signal_2086, signal_1190}), .c ({signal_2812, signal_1472}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1445 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2086, signal_1190}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1446 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2097, signal_1964}), .c ({signal_2140, signal_1189}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1447 ( .a ({signal_2813, signal_1191}), .b ({signal_2087, signal_1192}), .c ({signal_2844, signal_1473}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1448 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2087, signal_1192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1449 ( .a ({signal_2092, signal_1203}), .b ({signal_2143, signal_1965}), .c ({signal_2813, signal_1191}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1450 ( .a ({signal_2814, signal_1193}), .b ({signal_2088, signal_1194}), .c ({signal_2845, signal_1474}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1451 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2088, signal_1194}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1452 ( .a ({signal_2093, signal_1202}), .b ({signal_2144, signal_1966}), .c ({signal_2814, signal_1193}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1453 ( .a ({signal_2141, signal_1195}), .b ({signal_2089, signal_1196}), .c ({signal_2815, signal_1475}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1454 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2089, signal_1196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1455 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2098, signal_1967}), .c ({signal_2141, signal_1195}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1456 ( .a ({signal_2816, signal_1197}), .b ({signal_2090, signal_1198}), .c ({signal_2846, signal_1476}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1457 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2090, signal_1198}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1458 ( .a ({signal_2094, signal_1201}), .b ({signal_2145, signal_1968}), .c ({signal_2816, signal_1197}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1459 ( .a ({signal_2142, signal_1199}), .b ({signal_2091, signal_1200}), .c ({signal_2817, signal_1477}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1460 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2091, signal_1200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1461 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2099, signal_1969}), .c ({signal_2142, signal_1199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1462 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2092, signal_1203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1463 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2093, signal_1202}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1464 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2094, signal_1201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1465 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2095, signal_1962}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1466 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2096, signal_1963}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1467 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2097, signal_1964}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1468 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2100, signal_1970}), .c ({signal_2143, signal_1965}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1469 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2101, signal_1971}), .c ({signal_2144, signal_1966}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1470 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2098, signal_1967}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1471 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2102, signal_1973}), .c ({signal_2145, signal_1968}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1472 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2099, signal_1969}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1473 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2100, signal_1970}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1474 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2101, signal_1971}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1475 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2102, signal_1973}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1476 ( .a ({signal_2146, signal_1204}), .b ({signal_2103, signal_1205}), .c ({signal_2818, signal_1478}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1477 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2103, signal_1205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1478 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2114, signal_1974}), .c ({signal_2146, signal_1204}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1479 ( .a ({signal_2147, signal_1206}), .b ({signal_2104, signal_1207}), .c ({signal_2819, signal_1479}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1480 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2104, signal_1207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1481 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2115, signal_1975}), .c ({signal_2147, signal_1206}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1482 ( .a ({signal_2148, signal_1208}), .b ({signal_2105, signal_1209}), .c ({signal_2820, signal_1480}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1483 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2105, signal_1209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1484 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2116, signal_1976}), .c ({signal_2148, signal_1208}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1485 ( .a ({signal_2821, signal_1210}), .b ({signal_2106, signal_1211}), .c ({signal_2847, signal_1481}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1486 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2106, signal_1211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1487 ( .a ({signal_2111, signal_1222}), .b ({signal_2151, signal_1977}), .c ({signal_2821, signal_1210}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1488 ( .a ({signal_2822, signal_1212}), .b ({signal_2107, signal_1213}), .c ({signal_2848, signal_1482}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1489 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2107, signal_1213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1490 ( .a ({signal_2112, signal_1221}), .b ({signal_2152, signal_1978}), .c ({signal_2822, signal_1212}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1491 ( .a ({signal_2149, signal_1214}), .b ({signal_2108, signal_1215}), .c ({signal_2823, signal_1483}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1492 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2108, signal_1215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1493 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2117, signal_1979}), .c ({signal_2149, signal_1214}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1494 ( .a ({signal_2824, signal_1216}), .b ({signal_2109, signal_1217}), .c ({signal_2849, signal_1484}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1495 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2109, signal_1217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1496 ( .a ({signal_2113, signal_1220}), .b ({signal_2153, signal_1980}), .c ({signal_2824, signal_1216}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1497 ( .a ({signal_2150, signal_1218}), .b ({signal_2110, signal_1219}), .c ({signal_2825, signal_1485}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1498 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2110, signal_1219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1499 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2118, signal_1981}), .c ({signal_2150, signal_1218}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1500 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2111, signal_1222}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1501 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2112, signal_1221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1502 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2113, signal_1220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1503 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2114, signal_1974}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1504 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2115, signal_1975}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1505 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2116, signal_1976}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1506 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2119, signal_1225}), .c ({signal_2151, signal_1977}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1507 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2120, signal_1224}), .c ({signal_2152, signal_1978}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1508 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2117, signal_1979}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1509 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2121, signal_1223}), .c ({signal_2153, signal_1980}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1510 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2118, signal_1981}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1511 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2119, signal_1225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1512 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2120, signal_1224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1513 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2121, signal_1223}) ) ;
    NOR2_X1 cell_1514 ( .A1 (signal_1255), .A2 (signal_1226), .ZN (signal_1494) ) ;
    NOR2_X1 cell_1515 ( .A1 (signal_1257), .A2 (signal_1226), .ZN (signal_1495) ) ;
    AND2_X1 cell_1516 ( .A1 (signal_1273), .A2 (signal_397), .ZN (signal_1496) ) ;
    AND2_X1 cell_1517 ( .A1 (signal_1272), .A2 (signal_397), .ZN (signal_1497) ) ;
    NOR2_X1 cell_1518 ( .A1 (signal_1261), .A2 (signal_1226), .ZN (signal_1498) ) ;
    NOR2_X1 cell_1519 ( .A1 (signal_1263), .A2 (signal_1226), .ZN (signal_1499) ) ;
    NOR2_X1 cell_1520 ( .A1 (signal_1265), .A2 (signal_1226), .ZN (signal_1500) ) ;
    NOR2_X1 cell_1521 ( .A1 (signal_1267), .A2 (signal_1226), .ZN (signal_1501) ) ;
    INV_X1 cell_1522 ( .A (signal_397), .ZN (signal_1226) ) ;
    NAND2_X1 cell_1523 ( .A1 (signal_1227), .A2 (signal_1228), .ZN (signal_401) ) ;
    NOR2_X1 cell_1524 ( .A1 (signal_1229), .A2 (signal_1230), .ZN (signal_1228) ) ;
    NAND2_X1 cell_1525 ( .A1 (signal_1231), .A2 (signal_1232), .ZN (signal_1230) ) ;
    NOR2_X1 cell_1526 ( .A1 (signal_1269), .A2 (signal_1261), .ZN (signal_1232) ) ;
    NOR2_X1 cell_1527 ( .A1 (signal_1274), .A2 (signal_1267), .ZN (signal_1231) ) ;
    NAND2_X1 cell_1528 ( .A1 (signal_1270), .A2 (signal_1254), .ZN (signal_1229) ) ;
    NOR2_X1 cell_1529 ( .A1 (signal_1272), .A2 (signal_1273), .ZN (signal_1227) ) ;
    NAND2_X1 cell_1530 ( .A1 (signal_393), .A2 (signal_1233), .ZN (signal_1275) ) ;
    MUX2_X1 cell_1531 ( .S (signal_1253), .A (signal_1255), .B (signal_1267), .Z (signal_1233) ) ;
    NAND2_X1 cell_1532 ( .A1 (signal_1234), .A2 (signal_1235), .ZN (signal_1266) ) ;
    NAND2_X1 cell_1533 ( .A1 (signal_1236), .A2 (signal_1269), .ZN (signal_1235) ) ;
    NAND2_X1 cell_1534 ( .A1 (signal_1237), .A2 (signal_1238), .ZN (signal_1234) ) ;
    XOR2_X1 cell_1535 ( .A (signal_1268), .B (signal_1254), .Z (signal_1237) ) ;
    NAND2_X1 cell_1536 ( .A1 (signal_393), .A2 (signal_1239), .ZN (signal_1264) ) ;
    MUX2_X1 cell_1537 ( .S (signal_1253), .A (signal_1265), .B (signal_1263), .Z (signal_1239) ) ;
    NAND2_X1 cell_1538 ( .A1 (signal_393), .A2 (signal_1240), .ZN (signal_1262) ) ;
    MUX2_X1 cell_1539 ( .S (signal_1253), .A (signal_1241), .B (signal_1261), .Z (signal_1240) ) ;
    XNOR2_X1 cell_1540 ( .A (signal_1254), .B (signal_1270), .ZN (signal_1241) ) ;
    NAND2_X1 cell_1541 ( .A1 (signal_1242), .A2 (signal_1243), .ZN (signal_1260) ) ;
    NAND2_X1 cell_1542 ( .A1 (signal_1272), .A2 (signal_1236), .ZN (signal_1243) ) ;
    NAND2_X1 cell_1543 ( .A1 (signal_1244), .A2 (signal_1238), .ZN (signal_1242) ) ;
    XOR2_X1 cell_1544 ( .A (signal_1261), .B (signal_1255), .Z (signal_1244) ) ;
    NAND2_X1 cell_1545 ( .A1 (signal_1245), .A2 (signal_1246), .ZN (signal_1259) ) ;
    NAND2_X1 cell_1546 ( .A1 (signal_1272), .A2 (signal_1238), .ZN (signal_1246) ) ;
    NAND2_X1 cell_1547 ( .A1 (signal_1273), .A2 (signal_1236), .ZN (signal_1245) ) ;
    NAND2_X1 cell_1548 ( .A1 (signal_1247), .A2 (signal_1248), .ZN (signal_1258) ) ;
    NAND2_X1 cell_1549 ( .A1 (signal_1273), .A2 (signal_1238), .ZN (signal_1248) ) ;
    NOR2_X1 cell_1550 ( .A1 (signal_1253), .A2 (signal_1252), .ZN (signal_1238) ) ;
    NAND2_X1 cell_1551 ( .A1 (signal_1274), .A2 (signal_1236), .ZN (signal_1247) ) ;
    NOR2_X1 cell_1552 ( .A1 (signal_395), .A2 (signal_1252), .ZN (signal_1236) ) ;
    NAND2_X1 cell_1553 ( .A1 (signal_393), .A2 (signal_1249), .ZN (signal_1256) ) ;
    MUX2_X1 cell_1554 ( .S (signal_1253), .A (signal_1257), .B (signal_1255), .Z (signal_1249) ) ;
    NAND2_X1 cell_1555 ( .A1 (signal_1272), .A2 (signal_1270), .ZN (signal_1251) ) ;
    NAND2_X1 cell_1556 ( .A1 (signal_1269), .A2 (signal_1273), .ZN (signal_1250) ) ;
    INV_X1 cell_1557 ( .A (signal_393), .ZN (signal_1252) ) ;
    INV_X1 cell_1558 ( .A (signal_395), .ZN (signal_1253) ) ;
    NOR2_X1 cell_1559 ( .A1 (signal_1250), .A2 (signal_1251), .ZN (signal_399) ) ;
    INV_X1 cell_1560 ( .A (signal_1268), .ZN (signal_1267) ) ;
    INV_X1 cell_1562 ( .A (signal_1269), .ZN (signal_1265) ) ;
    INV_X1 cell_1564 ( .A (signal_1270), .ZN (signal_1263) ) ;
    INV_X1 cell_1566 ( .A (signal_1271), .ZN (signal_1261) ) ;
    INV_X1 cell_1572 ( .A (signal_1274), .ZN (signal_1257) ) ;
    INV_X1 cell_1574 ( .A (signal_1254), .ZN (signal_1255) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1576 ( .s (signal_394), .b ({signal_1984, signal_1413}), .a ({signal_2563, signal_1509}), .c ({signal_2826, signal_1517}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1577 ( .s (signal_394), .b ({signal_1987, signal_1412}), .a ({signal_2566, signal_1508}), .c ({signal_2827, signal_1516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1578 ( .s (signal_394), .b ({signal_1990, signal_1411}), .a ({signal_2569, signal_1507}), .c ({signal_2828, signal_1515}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1579 ( .s (signal_394), .b ({signal_1993, signal_1410}), .a ({signal_2572, signal_1506}), .c ({signal_2829, signal_1514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1580 ( .s (signal_394), .b ({signal_1996, signal_1409}), .a ({signal_2575, signal_1505}), .c ({signal_2830, signal_1513}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1581 ( .s (signal_394), .b ({signal_1999, signal_1408}), .a ({signal_2578, signal_1504}), .c ({signal_2831, signal_1512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1582 ( .s (signal_394), .b ({signal_2002, signal_1407}), .a ({signal_2581, signal_1503}), .c ({signal_2832, signal_1511}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1583 ( .s (signal_394), .b ({signal_2005, signal_1406}), .a ({signal_2584, signal_1502}), .c ({signal_2833, signal_1510}) ) ;
    INV_X1 cell_1712 ( .A (signal_393), .ZN (signal_402) ) ;
    ClockGatingController #(3) cell_1715 ( .clk (clk), .rst (start), .GatedClk (signal_3422), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_56 ( .s (signal_399), .b ({signal_2997, signal_1405}), .a ({signal_1984, signal_1413}), .c ({signal_2998, signal_1421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_57 ( .s (signal_399), .b ({signal_2996, signal_1404}), .a ({signal_1987, signal_1412}), .c ({signal_2999, signal_1420}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_58 ( .s (signal_399), .b ({signal_2995, signal_1403}), .a ({signal_1990, signal_1411}), .c ({signal_3000, signal_1419}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_59 ( .s (signal_399), .b ({signal_2994, signal_1402}), .a ({signal_1993, signal_1410}), .c ({signal_3001, signal_1418}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_60 ( .s (signal_399), .b ({signal_2993, signal_1401}), .a ({signal_1996, signal_1409}), .c ({signal_3002, signal_1417}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_61 ( .s (signal_399), .b ({signal_2992, signal_1400}), .a ({signal_1999, signal_1408}), .c ({signal_3003, signal_1416}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_62 ( .s (signal_399), .b ({signal_2991, signal_1399}), .a ({signal_2002, signal_1407}), .c ({signal_3004, signal_1415}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_63 ( .s (signal_399), .b ({signal_2990, signal_1398}), .a ({signal_2005, signal_1406}), .c ({signal_3005, signal_1414}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_445 ( .s (signal_464), .b ({signal_3247, signal_1557}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_3286, signal_705}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_448 ( .s (signal_464), .b ({signal_3249, signal_1556}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_3287, signal_707}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_451 ( .s (signal_464), .b ({signal_3251, signal_1555}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({signal_3288, signal_709}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_454 ( .s (signal_464), .b ({signal_3253, signal_1554}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({signal_3289, signal_711}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_457 ( .s (signal_464), .b ({signal_3255, signal_1553}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_3290, signal_713}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_460 ( .s (signal_464), .b ({signal_3257, signal_1552}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_3291, signal_715}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_463 ( .s (signal_464), .b ({signal_3259, signal_1551}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_3292, signal_717}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_466 ( .s (signal_464), .b ({signal_3261, signal_1550}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_3293, signal_719}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_613 ( .s (signal_455), .b ({signal_2998, signal_1421}), .a ({signal_2850, signal_1453}), .c ({signal_3086, signal_1525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_614 ( .s (signal_455), .b ({signal_2999, signal_1420}), .a ({signal_2851, signal_1452}), .c ({signal_3087, signal_1524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_615 ( .s (signal_455), .b ({signal_3000, signal_1419}), .a ({signal_2834, signal_1451}), .c ({signal_3088, signal_1523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_616 ( .s (signal_455), .b ({signal_3001, signal_1418}), .a ({signal_2852, signal_1450}), .c ({signal_3089, signal_1522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_617 ( .s (signal_455), .b ({signal_3002, signal_1417}), .a ({signal_2853, signal_1449}), .c ({signal_3090, signal_1521}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_618 ( .s (signal_455), .b ({signal_3003, signal_1416}), .a ({signal_2835, signal_1448}), .c ({signal_3091, signal_1520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_619 ( .s (signal_455), .b ({signal_3004, signal_1415}), .a ({signal_2836, signal_1447}), .c ({signal_3092, signal_1519}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_620 ( .s (signal_455), .b ({signal_3005, signal_1414}), .a ({signal_2837, signal_1446}), .c ({signal_3093, signal_1518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_621 ( .s (signal_452), .b ({plaintext_s1[0], plaintext_s0[0]}), .a ({signal_3086, signal_1525}), .c ({signal_3247, signal_1557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_622 ( .s (signal_452), .b ({plaintext_s1[1], plaintext_s0[1]}), .a ({signal_3087, signal_1524}), .c ({signal_3249, signal_1556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_623 ( .s (signal_452), .b ({plaintext_s1[2], plaintext_s0[2]}), .a ({signal_3088, signal_1523}), .c ({signal_3251, signal_1555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_624 ( .s (signal_452), .b ({plaintext_s1[3], plaintext_s0[3]}), .a ({signal_3089, signal_1522}), .c ({signal_3253, signal_1554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_625 ( .s (signal_452), .b ({plaintext_s1[4], plaintext_s0[4]}), .a ({signal_3090, signal_1521}), .c ({signal_3255, signal_1553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_626 ( .s (signal_452), .b ({plaintext_s1[5], plaintext_s0[5]}), .a ({signal_3091, signal_1520}), .c ({signal_3257, signal_1552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_627 ( .s (signal_452), .b ({plaintext_s1[6], plaintext_s0[6]}), .a ({signal_3092, signal_1519}), .c ({signal_3259, signal_1551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_628 ( .s (signal_452), .b ({plaintext_s1[7], plaintext_s0[7]}), .a ({signal_3093, signal_1518}), .c ({signal_3261, signal_1550}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_672 ( .a ({signal_3030, signal_724}), .b ({signal_2004, signal_1486}), .c ({signal_3094, signal_1750}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_673 ( .a ({1'b0, signal_1494}), .b ({signal_2990, signal_1398}), .c ({signal_3030, signal_724}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_674 ( .a ({signal_3031, signal_725}), .b ({signal_2001, signal_1487}), .c ({signal_3095, signal_1751}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_675 ( .a ({1'b0, signal_1495}), .b ({signal_2991, signal_1399}), .c ({signal_3031, signal_725}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_676 ( .a ({signal_3032, signal_726}), .b ({signal_1998, signal_1488}), .c ({signal_3096, signal_1752}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_677 ( .a ({1'b0, signal_1496}), .b ({signal_2992, signal_1400}), .c ({signal_3032, signal_726}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_678 ( .a ({signal_3033, signal_727}), .b ({signal_1995, signal_1489}), .c ({signal_3097, signal_1753}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_679 ( .a ({1'b0, signal_1497}), .b ({signal_2993, signal_1401}), .c ({signal_3033, signal_727}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_680 ( .a ({signal_3034, signal_728}), .b ({signal_1992, signal_1490}), .c ({signal_3098, signal_1754}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_681 ( .a ({1'b0, signal_1498}), .b ({signal_2994, signal_1402}), .c ({signal_3034, signal_728}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_682 ( .a ({signal_3035, signal_729}), .b ({signal_1989, signal_1491}), .c ({signal_3099, signal_1755}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_683 ( .a ({1'b0, signal_1499}), .b ({signal_2995, signal_1403}), .c ({signal_3035, signal_729}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_684 ( .a ({signal_3036, signal_730}), .b ({signal_1986, signal_1492}), .c ({signal_3100, signal_1756}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_685 ( .a ({1'b0, signal_1500}), .b ({signal_2996, signal_1404}), .c ({signal_3036, signal_730}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_686 ( .a ({signal_3037, signal_731}), .b ({signal_1983, signal_1493}), .c ({signal_3101, signal_1757}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_687 ( .a ({1'b0, signal_1501}), .b ({signal_2997, signal_1405}), .c ({signal_3037, signal_731}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1098 ( .s (signal_756), .b ({signal_2683, signal_1749}), .a ({signal_3262, signal_1055}), .c ({signal_3374, signal_1054}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1099 ( .s (signal_748), .b ({signal_2708, signal_1765}), .a ({signal_3101, signal_1757}), .c ({signal_3262, signal_1055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1102 ( .s (signal_756), .b ({signal_2686, signal_1748}), .a ({signal_3263, signal_1058}), .c ({signal_3375, signal_1057}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1103 ( .s (signal_748), .b ({signal_2711, signal_1764}), .a ({signal_3100, signal_1756}), .c ({signal_3263, signal_1058}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1106 ( .s (signal_756), .b ({signal_2689, signal_1747}), .a ({signal_3264, signal_1061}), .c ({signal_3376, signal_1060}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1107 ( .s (signal_748), .b ({signal_2714, signal_1763}), .a ({signal_3099, signal_1755}), .c ({signal_3264, signal_1061}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1110 ( .s (signal_756), .b ({signal_2692, signal_1746}), .a ({signal_3265, signal_1064}), .c ({signal_3377, signal_1063}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1111 ( .s (signal_748), .b ({signal_2717, signal_1762}), .a ({signal_3098, signal_1754}), .c ({signal_3265, signal_1064}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1114 ( .s (signal_756), .b ({signal_2695, signal_1745}), .a ({signal_3266, signal_1067}), .c ({signal_3378, signal_1066}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1115 ( .s (signal_748), .b ({signal_2720, signal_1761}), .a ({signal_3097, signal_1753}), .c ({signal_3266, signal_1067}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1118 ( .s (signal_756), .b ({signal_2698, signal_1744}), .a ({signal_3267, signal_1070}), .c ({signal_3379, signal_1069}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1119 ( .s (signal_748), .b ({signal_2723, signal_1760}), .a ({signal_3096, signal_1752}), .c ({signal_3267, signal_1070}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1122 ( .s (signal_756), .b ({signal_2701, signal_1743}), .a ({signal_3268, signal_1073}), .c ({signal_3380, signal_1072}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1123 ( .s (signal_748), .b ({signal_2726, signal_1759}), .a ({signal_3095, signal_1751}), .c ({signal_3268, signal_1073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1126 ( .s (signal_756), .b ({signal_2704, signal_1742}), .a ({signal_3269, signal_1076}), .c ({signal_3381, signal_1075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1127 ( .s (signal_748), .b ({signal_2729, signal_1758}), .a ({signal_3094, signal_1750}), .c ({signal_3269, signal_1076}) ) ;
    AES_step2_ANF #(.low_latency(0), .pipeline(0)) cell_1714 ( .in0 ({signal_1517, signal_1516, signal_1515, signal_1514, signal_1513, signal_1512, signal_1511, signal_1510}), .in1 ({signal_2826, signal_2827, signal_2828, signal_2829, signal_2830, signal_2831, signal_2832, signal_2833}), .clk (clk), .r ({Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_1405, signal_1404, signal_1403, signal_1402, signal_1401, signal_1400, signal_1399, signal_1398}), .out1 ({signal_2997, signal_2996, signal_2995, signal_2994, signal_2993, signal_2992, signal_2991, signal_2990}) ) ;

    /* register cells */
    DFF_X1 cell_33 ( .CK (signal_3422), .D (signal_429), .Q (signal_425), .QN () ) ;
    DFF_X1 cell_36 ( .CK (signal_3422), .D (signal_431), .Q (signal_426), .QN () ) ;
    DFF_X1 cell_39 ( .CK (signal_3422), .D (signal_433), .Q (signal_427), .QN () ) ;
    DFF_X1 cell_42 ( .CK (signal_3422), .D (signal_435), .Q (signal_428), .QN () ) ;
    DFF_X1 cell_45 ( .CK (signal_3422), .D (signal_437), .Q (signal_424), .QN () ) ;
    DFF_X1 cell_48 ( .CK (signal_3422), .D (signal_439), .Q (signal_421), .QN () ) ;
    DFF_X1 cell_51 ( .CK (signal_3422), .D (signal_441), .Q (signal_420), .QN () ) ;
    DFF_X1 cell_53 ( .CK (signal_3422), .D (signal_419), .Q (signal_418), .QN () ) ;
    DFF_X1 cell_55 ( .CK (signal_3422), .D (signal_395), .Q (signal_397), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_87 ( .clk (signal_3422), .D ({signal_3126, signal_465}), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_90 ( .clk (signal_3422), .D ({signal_3127, signal_467}), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_93 ( .clk (signal_3422), .D ({signal_3128, signal_469}), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_96 ( .clk (signal_3422), .D ({signal_3129, signal_471}), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_99 ( .clk (signal_3422), .D ({signal_3130, signal_473}), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_102 ( .clk (signal_3422), .D ({signal_3131, signal_475}), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_105 ( .clk (signal_3422), .D ({signal_3132, signal_477}), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_108 ( .clk (signal_3422), .D ({signal_3133, signal_479}), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_111 ( .clk (signal_3422), .D ({signal_3134, signal_481}), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_114 ( .clk (signal_3422), .D ({signal_3135, signal_483}), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_117 ( .clk (signal_3422), .D ({signal_3136, signal_485}), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_120 ( .clk (signal_3422), .D ({signal_3137, signal_487}), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_123 ( .clk (signal_3422), .D ({signal_3138, signal_489}), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_126 ( .clk (signal_3422), .D ({signal_3139, signal_491}), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_129 ( .clk (signal_3422), .D ({signal_3140, signal_493}), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_132 ( .clk (signal_3422), .D ({signal_3141, signal_495}), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_135 ( .clk (signal_3422), .D ({signal_3142, signal_497}), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_138 ( .clk (signal_3422), .D ({signal_3143, signal_499}), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_141 ( .clk (signal_3422), .D ({signal_3144, signal_501}), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_144 ( .clk (signal_3422), .D ({signal_3145, signal_503}), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_147 ( .clk (signal_3422), .D ({signal_3146, signal_505}), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_150 ( .clk (signal_3422), .D ({signal_3147, signal_507}), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_153 ( .clk (signal_3422), .D ({signal_3148, signal_509}), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_156 ( .clk (signal_3422), .D ({signal_3149, signal_511}), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_159 ( .clk (signal_3422), .D ({signal_3150, signal_513}), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_162 ( .clk (signal_3422), .D ({signal_3151, signal_515}), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_165 ( .clk (signal_3422), .D ({signal_3152, signal_517}), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_168 ( .clk (signal_3422), .D ({signal_3153, signal_519}), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_171 ( .clk (signal_3422), .D ({signal_3154, signal_521}), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_174 ( .clk (signal_3422), .D ({signal_3155, signal_523}), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_177 ( .clk (signal_3422), .D ({signal_3156, signal_525}), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_180 ( .clk (signal_3422), .D ({signal_3157, signal_527}), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_183 ( .clk (signal_3422), .D ({signal_3158, signal_529}), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_186 ( .clk (signal_3422), .D ({signal_3159, signal_531}), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_189 ( .clk (signal_3422), .D ({signal_3160, signal_533}), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_192 ( .clk (signal_3422), .D ({signal_3161, signal_535}), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_195 ( .clk (signal_3422), .D ({signal_3162, signal_537}), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_198 ( .clk (signal_3422), .D ({signal_3163, signal_539}), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_201 ( .clk (signal_3422), .D ({signal_3164, signal_541}), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_204 ( .clk (signal_3422), .D ({signal_3165, signal_543}), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_207 ( .clk (signal_3422), .D ({signal_3166, signal_545}), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_210 ( .clk (signal_3422), .D ({signal_3167, signal_547}), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_213 ( .clk (signal_3422), .D ({signal_3168, signal_549}), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_216 ( .clk (signal_3422), .D ({signal_3169, signal_551}), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_219 ( .clk (signal_3422), .D ({signal_3170, signal_553}), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_222 ( .clk (signal_3422), .D ({signal_3171, signal_555}), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_225 ( .clk (signal_3422), .D ({signal_3172, signal_557}), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_228 ( .clk (signal_3422), .D ({signal_3173, signal_559}), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_231 ( .clk (signal_3422), .D ({signal_3174, signal_561}), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_234 ( .clk (signal_3422), .D ({signal_3175, signal_563}), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_237 ( .clk (signal_3422), .D ({signal_3176, signal_565}), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_240 ( .clk (signal_3422), .D ({signal_3177, signal_567}), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_243 ( .clk (signal_3422), .D ({signal_3178, signal_569}), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_246 ( .clk (signal_3422), .D ({signal_3179, signal_571}), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_249 ( .clk (signal_3422), .D ({signal_3180, signal_573}), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_252 ( .clk (signal_3422), .D ({signal_3181, signal_575}), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_255 ( .clk (signal_3422), .D ({signal_3182, signal_577}), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_258 ( .clk (signal_3422), .D ({signal_3183, signal_579}), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_261 ( .clk (signal_3422), .D ({signal_3184, signal_581}), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_264 ( .clk (signal_3422), .D ({signal_3185, signal_583}), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_267 ( .clk (signal_3422), .D ({signal_3186, signal_585}), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_270 ( .clk (signal_3422), .D ({signal_3187, signal_587}), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_273 ( .clk (signal_3422), .D ({signal_3188, signal_589}), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_276 ( .clk (signal_3422), .D ({signal_3189, signal_591}), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_279 ( .clk (signal_3422), .D ({signal_3190, signal_593}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_282 ( .clk (signal_3422), .D ({signal_3191, signal_595}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_285 ( .clk (signal_3422), .D ({signal_3192, signal_597}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_288 ( .clk (signal_3422), .D ({signal_3193, signal_599}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_291 ( .clk (signal_3422), .D ({signal_3194, signal_601}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_294 ( .clk (signal_3422), .D ({signal_3195, signal_603}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_297 ( .clk (signal_3422), .D ({signal_3196, signal_605}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_300 ( .clk (signal_3422), .D ({signal_3197, signal_607}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_303 ( .clk (signal_3422), .D ({signal_3198, signal_609}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_306 ( .clk (signal_3422), .D ({signal_3199, signal_611}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_309 ( .clk (signal_3422), .D ({signal_3200, signal_613}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_312 ( .clk (signal_3422), .D ({signal_3201, signal_615}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_315 ( .clk (signal_3422), .D ({signal_3202, signal_617}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_318 ( .clk (signal_3422), .D ({signal_3203, signal_619}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_321 ( .clk (signal_3422), .D ({signal_3204, signal_621}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_324 ( .clk (signal_3422), .D ({signal_3205, signal_623}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_327 ( .clk (signal_3422), .D ({signal_3206, signal_625}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_330 ( .clk (signal_3422), .D ({signal_3207, signal_627}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_333 ( .clk (signal_3422), .D ({signal_3208, signal_629}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_336 ( .clk (signal_3422), .D ({signal_3209, signal_631}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_339 ( .clk (signal_3422), .D ({signal_3210, signal_633}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_342 ( .clk (signal_3422), .D ({signal_3211, signal_635}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_345 ( .clk (signal_3422), .D ({signal_3212, signal_637}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_348 ( .clk (signal_3422), .D ({signal_3213, signal_639}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_351 ( .clk (signal_3422), .D ({signal_3214, signal_641}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_354 ( .clk (signal_3422), .D ({signal_3215, signal_643}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_357 ( .clk (signal_3422), .D ({signal_3216, signal_645}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_360 ( .clk (signal_3422), .D ({signal_3217, signal_647}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_363 ( .clk (signal_3422), .D ({signal_3218, signal_649}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_366 ( .clk (signal_3422), .D ({signal_3219, signal_651}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_369 ( .clk (signal_3422), .D ({signal_3220, signal_653}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_372 ( .clk (signal_3422), .D ({signal_3221, signal_655}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_375 ( .clk (signal_3422), .D ({signal_3222, signal_657}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_378 ( .clk (signal_3422), .D ({signal_3223, signal_659}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_381 ( .clk (signal_3422), .D ({signal_3224, signal_661}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_384 ( .clk (signal_3422), .D ({signal_3225, signal_663}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_387 ( .clk (signal_3422), .D ({signal_3226, signal_665}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_390 ( .clk (signal_3422), .D ({signal_3227, signal_667}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_393 ( .clk (signal_3422), .D ({signal_3228, signal_669}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_396 ( .clk (signal_3422), .D ({signal_3229, signal_671}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_399 ( .clk (signal_3422), .D ({signal_3230, signal_673}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_402 ( .clk (signal_3422), .D ({signal_3231, signal_675}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_405 ( .clk (signal_3422), .D ({signal_3232, signal_677}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_408 ( .clk (signal_3422), .D ({signal_3233, signal_679}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_411 ( .clk (signal_3422), .D ({signal_3234, signal_681}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_414 ( .clk (signal_3422), .D ({signal_3235, signal_683}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_417 ( .clk (signal_3422), .D ({signal_3236, signal_685}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_420 ( .clk (signal_3422), .D ({signal_3237, signal_687}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_423 ( .clk (signal_3422), .D ({signal_3238, signal_689}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_426 ( .clk (signal_3422), .D ({signal_3239, signal_691}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_429 ( .clk (signal_3422), .D ({signal_3240, signal_693}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_432 ( .clk (signal_3422), .D ({signal_3241, signal_695}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_435 ( .clk (signal_3422), .D ({signal_3242, signal_697}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_438 ( .clk (signal_3422), .D ({signal_3243, signal_699}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_441 ( .clk (signal_3422), .D ({signal_3244, signal_701}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_444 ( .clk (signal_3422), .D ({signal_3245, signal_703}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_447 ( .clk (signal_3422), .D ({signal_3286, signal_705}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_450 ( .clk (signal_3422), .D ({signal_3287, signal_707}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_453 ( .clk (signal_3422), .D ({signal_3288, signal_709}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_456 ( .clk (signal_3422), .D ({signal_3289, signal_711}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_459 ( .clk (signal_3422), .D ({signal_3290, signal_713}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_462 ( .clk (signal_3422), .D ({signal_3291, signal_715}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_465 ( .clk (signal_3422), .D ({signal_3292, signal_717}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_468 ( .clk (signal_3422), .D ({signal_3293, signal_719}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_717 ( .clk (signal_3422), .D ({signal_3406, signal_766}), .Q ({signal_1983, signal_1493}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_721 ( .clk (signal_3422), .D ({signal_3407, signal_769}), .Q ({signal_1986, signal_1492}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_725 ( .clk (signal_3422), .D ({signal_3408, signal_772}), .Q ({signal_1989, signal_1491}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_729 ( .clk (signal_3422), .D ({signal_3409, signal_775}), .Q ({signal_1992, signal_1490}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_733 ( .clk (signal_3422), .D ({signal_3410, signal_778}), .Q ({signal_1995, signal_1489}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_737 ( .clk (signal_3422), .D ({signal_3411, signal_781}), .Q ({signal_1998, signal_1488}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_741 ( .clk (signal_3422), .D ({signal_3412, signal_784}), .Q ({signal_2001, signal_1487}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_745 ( .clk (signal_3422), .D ({signal_3413, signal_787}), .Q ({signal_2004, signal_1486}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_749 ( .clk (signal_3422), .D ({signal_3302, signal_790}), .Q ({signal_2020, signal_758}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_753 ( .clk (signal_3422), .D ({signal_3303, signal_793}), .Q ({signal_2018, signal_759}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_757 ( .clk (signal_3422), .D ({signal_3304, signal_796}), .Q ({signal_2016, signal_760}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_761 ( .clk (signal_3422), .D ({signal_3305, signal_799}), .Q ({signal_2014, signal_761}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_765 ( .clk (signal_3422), .D ({signal_3306, signal_802}), .Q ({signal_2012, signal_762}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_769 ( .clk (signal_3422), .D ({signal_3307, signal_805}), .Q ({signal_2010, signal_763}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_773 ( .clk (signal_3422), .D ({signal_3308, signal_808}), .Q ({signal_2008, signal_764}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_777 ( .clk (signal_3422), .D ({signal_3309, signal_811}), .Q ({signal_2006, signal_765}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_781 ( .clk (signal_3422), .D ({signal_3310, signal_814}), .Q ({signal_2443, signal_1909}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_785 ( .clk (signal_3422), .D ({signal_3311, signal_817}), .Q ({signal_2446, signal_1908}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_789 ( .clk (signal_3422), .D ({signal_3312, signal_820}), .Q ({signal_2449, signal_1907}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_793 ( .clk (signal_3422), .D ({signal_3313, signal_823}), .Q ({signal_2452, signal_1906}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_797 ( .clk (signal_3422), .D ({signal_3314, signal_826}), .Q ({signal_2455, signal_1905}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_801 ( .clk (signal_3422), .D ({signal_3315, signal_829}), .Q ({signal_2458, signal_1904}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_805 ( .clk (signal_3422), .D ({signal_3316, signal_832}), .Q ({signal_2461, signal_1903}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_809 ( .clk (signal_3422), .D ({signal_3317, signal_835}), .Q ({signal_2464, signal_1902}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_813 ( .clk (signal_3422), .D ({signal_3318, signal_838}), .Q ({signal_2467, signal_1893}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_817 ( .clk (signal_3422), .D ({signal_3319, signal_841}), .Q ({signal_2470, signal_1892}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_821 ( .clk (signal_3422), .D ({signal_3320, signal_844}), .Q ({signal_2473, signal_1891}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_825 ( .clk (signal_3422), .D ({signal_3321, signal_847}), .Q ({signal_2476, signal_1890}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_829 ( .clk (signal_3422), .D ({signal_3322, signal_850}), .Q ({signal_2479, signal_1889}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_833 ( .clk (signal_3422), .D ({signal_3323, signal_853}), .Q ({signal_2482, signal_1888}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_837 ( .clk (signal_3422), .D ({signal_3324, signal_856}), .Q ({signal_2485, signal_1887}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_841 ( .clk (signal_3422), .D ({signal_3325, signal_859}), .Q ({signal_2488, signal_1886}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_845 ( .clk (signal_3422), .D ({signal_3326, signal_862}), .Q ({signal_2491, signal_1877}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_849 ( .clk (signal_3422), .D ({signal_3327, signal_865}), .Q ({signal_2494, signal_1876}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_853 ( .clk (signal_3422), .D ({signal_3328, signal_868}), .Q ({signal_2497, signal_1875}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_857 ( .clk (signal_3422), .D ({signal_3329, signal_871}), .Q ({signal_2500, signal_1874}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_861 ( .clk (signal_3422), .D ({signal_3330, signal_874}), .Q ({signal_2503, signal_1873}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_865 ( .clk (signal_3422), .D ({signal_3331, signal_877}), .Q ({signal_2506, signal_1872}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_869 ( .clk (signal_3422), .D ({signal_3332, signal_880}), .Q ({signal_2509, signal_1871}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_873 ( .clk (signal_3422), .D ({signal_3333, signal_883}), .Q ({signal_2512, signal_1870}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_877 ( .clk (signal_3422), .D ({signal_3334, signal_886}), .Q ({signal_2515, signal_1861}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_881 ( .clk (signal_3422), .D ({signal_3335, signal_889}), .Q ({signal_2518, signal_1860}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_885 ( .clk (signal_3422), .D ({signal_3336, signal_892}), .Q ({signal_2521, signal_1859}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_889 ( .clk (signal_3422), .D ({signal_3337, signal_895}), .Q ({signal_2524, signal_1858}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_893 ( .clk (signal_3422), .D ({signal_3338, signal_898}), .Q ({signal_2527, signal_1857}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_897 ( .clk (signal_3422), .D ({signal_3339, signal_901}), .Q ({signal_2530, signal_1856}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_901 ( .clk (signal_3422), .D ({signal_3340, signal_904}), .Q ({signal_2533, signal_1855}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_905 ( .clk (signal_3422), .D ({signal_3341, signal_907}), .Q ({signal_2536, signal_1854}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_909 ( .clk (signal_3422), .D ({signal_3102, signal_910}), .Q ({signal_2539, signal_1845}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_913 ( .clk (signal_3422), .D ({signal_3103, signal_913}), .Q ({signal_2542, signal_1844}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_917 ( .clk (signal_3422), .D ({signal_3104, signal_916}), .Q ({signal_2545, signal_1843}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_921 ( .clk (signal_3422), .D ({signal_3105, signal_919}), .Q ({signal_2548, signal_1842}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_925 ( .clk (signal_3422), .D ({signal_3106, signal_922}), .Q ({signal_2551, signal_1841}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_929 ( .clk (signal_3422), .D ({signal_3107, signal_925}), .Q ({signal_2554, signal_1840}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_933 ( .clk (signal_3422), .D ({signal_3108, signal_928}), .Q ({signal_2557, signal_1839}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_937 ( .clk (signal_3422), .D ({signal_3109, signal_931}), .Q ({signal_2560, signal_1838}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_941 ( .clk (signal_3422), .D ({signal_3110, signal_934}), .Q ({signal_2563, signal_1509}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_945 ( .clk (signal_3422), .D ({signal_3111, signal_937}), .Q ({signal_2566, signal_1508}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_949 ( .clk (signal_3422), .D ({signal_3112, signal_940}), .Q ({signal_2569, signal_1507}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_953 ( .clk (signal_3422), .D ({signal_3113, signal_943}), .Q ({signal_2572, signal_1506}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_957 ( .clk (signal_3422), .D ({signal_3114, signal_946}), .Q ({signal_2575, signal_1505}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_961 ( .clk (signal_3422), .D ({signal_3115, signal_949}), .Q ({signal_2578, signal_1504}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_965 ( .clk (signal_3422), .D ({signal_3116, signal_952}), .Q ({signal_2581, signal_1503}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_969 ( .clk (signal_3422), .D ({signal_3117, signal_955}), .Q ({signal_2584, signal_1502}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_973 ( .clk (signal_3422), .D ({signal_3342, signal_958}), .Q ({signal_2587, signal_1821}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_977 ( .clk (signal_3422), .D ({signal_3343, signal_961}), .Q ({signal_2590, signal_1820}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_981 ( .clk (signal_3422), .D ({signal_3344, signal_964}), .Q ({signal_2593, signal_1819}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_985 ( .clk (signal_3422), .D ({signal_3345, signal_967}), .Q ({signal_2596, signal_1818}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_989 ( .clk (signal_3422), .D ({signal_3346, signal_970}), .Q ({signal_2599, signal_1817}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_993 ( .clk (signal_3422), .D ({signal_3347, signal_973}), .Q ({signal_2602, signal_1816}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_997 ( .clk (signal_3422), .D ({signal_3348, signal_976}), .Q ({signal_2605, signal_1815}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1001 ( .clk (signal_3422), .D ({signal_3349, signal_979}), .Q ({signal_2608, signal_1814}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1005 ( .clk (signal_3422), .D ({signal_3350, signal_982}), .Q ({signal_2611, signal_1805}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1009 ( .clk (signal_3422), .D ({signal_3351, signal_985}), .Q ({signal_2614, signal_1804}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1013 ( .clk (signal_3422), .D ({signal_3352, signal_988}), .Q ({signal_2617, signal_1803}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1017 ( .clk (signal_3422), .D ({signal_3353, signal_991}), .Q ({signal_2620, signal_1802}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1021 ( .clk (signal_3422), .D ({signal_3354, signal_994}), .Q ({signal_2623, signal_1801}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1025 ( .clk (signal_3422), .D ({signal_3355, signal_997}), .Q ({signal_2626, signal_1800}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1029 ( .clk (signal_3422), .D ({signal_3356, signal_1000}), .Q ({signal_2629, signal_1799}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1033 ( .clk (signal_3422), .D ({signal_3357, signal_1003}), .Q ({signal_2632, signal_1798}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1037 ( .clk (signal_3422), .D ({signal_3358, signal_1006}), .Q ({signal_2635, signal_1789}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1041 ( .clk (signal_3422), .D ({signal_3359, signal_1009}), .Q ({signal_2638, signal_1788}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1045 ( .clk (signal_3422), .D ({signal_3360, signal_1012}), .Q ({signal_2641, signal_1787}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1049 ( .clk (signal_3422), .D ({signal_3361, signal_1015}), .Q ({signal_2644, signal_1786}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1053 ( .clk (signal_3422), .D ({signal_3362, signal_1018}), .Q ({signal_2647, signal_1785}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1057 ( .clk (signal_3422), .D ({signal_3363, signal_1021}), .Q ({signal_2650, signal_1784}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1061 ( .clk (signal_3422), .D ({signal_3364, signal_1024}), .Q ({signal_2653, signal_1783}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1065 ( .clk (signal_3422), .D ({signal_3365, signal_1027}), .Q ({signal_2656, signal_1782}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1069 ( .clk (signal_3422), .D ({signal_3366, signal_1030}), .Q ({signal_2659, signal_1773}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1073 ( .clk (signal_3422), .D ({signal_3367, signal_1033}), .Q ({signal_2662, signal_1772}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1077 ( .clk (signal_3422), .D ({signal_3368, signal_1036}), .Q ({signal_2665, signal_1771}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1081 ( .clk (signal_3422), .D ({signal_3369, signal_1039}), .Q ({signal_2668, signal_1770}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1085 ( .clk (signal_3422), .D ({signal_3370, signal_1042}), .Q ({signal_2671, signal_1769}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1089 ( .clk (signal_3422), .D ({signal_3371, signal_1045}), .Q ({signal_2674, signal_1768}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1093 ( .clk (signal_3422), .D ({signal_3372, signal_1048}), .Q ({signal_2677, signal_1767}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1097 ( .clk (signal_3422), .D ({signal_3373, signal_1051}), .Q ({signal_2680, signal_1766}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1101 ( .clk (signal_3422), .D ({signal_3374, signal_1054}), .Q ({signal_2683, signal_1749}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1105 ( .clk (signal_3422), .D ({signal_3375, signal_1057}), .Q ({signal_2686, signal_1748}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1109 ( .clk (signal_3422), .D ({signal_3376, signal_1060}), .Q ({signal_2689, signal_1747}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1113 ( .clk (signal_3422), .D ({signal_3377, signal_1063}), .Q ({signal_2692, signal_1746}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1117 ( .clk (signal_3422), .D ({signal_3378, signal_1066}), .Q ({signal_2695, signal_1745}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1121 ( .clk (signal_3422), .D ({signal_3379, signal_1069}), .Q ({signal_2698, signal_1744}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1125 ( .clk (signal_3422), .D ({signal_3380, signal_1072}), .Q ({signal_2701, signal_1743}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1129 ( .clk (signal_3422), .D ({signal_3381, signal_1075}), .Q ({signal_2704, signal_1742}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1133 ( .clk (signal_3422), .D ({signal_3382, signal_1078}), .Q ({signal_2707, signal_1733}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1137 ( .clk (signal_3422), .D ({signal_3383, signal_1081}), .Q ({signal_2710, signal_1732}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1141 ( .clk (signal_3422), .D ({signal_3384, signal_1084}), .Q ({signal_2713, signal_1731}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1145 ( .clk (signal_3422), .D ({signal_3385, signal_1087}), .Q ({signal_2716, signal_1730}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1149 ( .clk (signal_3422), .D ({signal_3386, signal_1090}), .Q ({signal_2719, signal_1729}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1153 ( .clk (signal_3422), .D ({signal_3387, signal_1093}), .Q ({signal_2722, signal_1728}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1157 ( .clk (signal_3422), .D ({signal_3388, signal_1096}), .Q ({signal_2725, signal_1727}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1161 ( .clk (signal_3422), .D ({signal_3389, signal_1099}), .Q ({signal_2728, signal_1726}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1165 ( .clk (signal_3422), .D ({signal_3390, signal_1102}), .Q ({signal_2731, signal_1717}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1169 ( .clk (signal_3422), .D ({signal_3391, signal_1105}), .Q ({signal_2734, signal_1716}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1173 ( .clk (signal_3422), .D ({signal_3392, signal_1108}), .Q ({signal_2737, signal_1715}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1177 ( .clk (signal_3422), .D ({signal_3393, signal_1111}), .Q ({signal_2740, signal_1714}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1181 ( .clk (signal_3422), .D ({signal_3394, signal_1114}), .Q ({signal_2743, signal_1713}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1185 ( .clk (signal_3422), .D ({signal_3395, signal_1117}), .Q ({signal_2746, signal_1712}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1189 ( .clk (signal_3422), .D ({signal_3396, signal_1120}), .Q ({signal_2749, signal_1711}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1193 ( .clk (signal_3422), .D ({signal_3397, signal_1123}), .Q ({signal_2752, signal_1710}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1197 ( .clk (signal_3422), .D ({signal_3398, signal_1126}), .Q ({signal_2755, signal_1701}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1201 ( .clk (signal_3422), .D ({signal_3399, signal_1129}), .Q ({signal_2758, signal_1700}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1205 ( .clk (signal_3422), .D ({signal_3400, signal_1132}), .Q ({signal_2761, signal_1699}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1209 ( .clk (signal_3422), .D ({signal_3401, signal_1135}), .Q ({signal_2764, signal_1698}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1213 ( .clk (signal_3422), .D ({signal_3402, signal_1138}), .Q ({signal_2767, signal_1697}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1217 ( .clk (signal_3422), .D ({signal_3403, signal_1141}), .Q ({signal_2770, signal_1696}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1221 ( .clk (signal_3422), .D ({signal_3404, signal_1144}), .Q ({signal_2773, signal_1695}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1225 ( .clk (signal_3422), .D ({signal_3405, signal_1147}), .Q ({signal_2776, signal_1694}) ) ;
    DFF_X1 cell_1561 ( .CK (signal_3422), .D (signal_1275), .Q (signal_1268), .QN () ) ;
    DFF_X1 cell_1563 ( .CK (signal_3422), .D (signal_1266), .Q (signal_1269), .QN () ) ;
    DFF_X1 cell_1565 ( .CK (signal_3422), .D (signal_1264), .Q (signal_1270), .QN () ) ;
    DFF_X1 cell_1567 ( .CK (signal_3422), .D (signal_1262), .Q (signal_1271), .QN () ) ;
    DFF_X1 cell_1569 ( .CK (signal_3422), .D (signal_1260), .Q (signal_1272), .QN () ) ;
    DFF_X1 cell_1571 ( .CK (signal_3422), .D (signal_1259), .Q (signal_1273), .QN () ) ;
    DFF_X1 cell_1573 ( .CK (signal_3422), .D (signal_1258), .Q (signal_1274), .QN () ) ;
    DFF_X1 cell_1575 ( .CK (signal_3422), .D (signal_1256), .Q (signal_1254), .QN () ) ;
    DFF_X1 cell_1713 ( .CK (signal_3422), .D (signal_403), .Q (signal_393), .QN () ) ;
endmodule
