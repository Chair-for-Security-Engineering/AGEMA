////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_round-based/AGEMA/AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d2 (plaintext_s0, key_s0, clk, reset, key_s1, key_s2, plaintext_s1, plaintext_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [4079:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_16933 ;
    wire new_AGEMA_signal_16934 ;
    wire new_AGEMA_signal_16935 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16939 ;
    wire new_AGEMA_signal_16940 ;
    wire new_AGEMA_signal_16941 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16945 ;
    wire new_AGEMA_signal_16946 ;
    wire new_AGEMA_signal_16947 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16951 ;
    wire new_AGEMA_signal_16952 ;
    wire new_AGEMA_signal_16953 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16957 ;
    wire new_AGEMA_signal_16958 ;
    wire new_AGEMA_signal_16959 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16963 ;
    wire new_AGEMA_signal_16964 ;
    wire new_AGEMA_signal_16965 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16969 ;
    wire new_AGEMA_signal_16970 ;
    wire new_AGEMA_signal_16971 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16975 ;
    wire new_AGEMA_signal_16976 ;
    wire new_AGEMA_signal_16977 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16981 ;
    wire new_AGEMA_signal_16982 ;
    wire new_AGEMA_signal_16983 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16987 ;
    wire new_AGEMA_signal_16988 ;
    wire new_AGEMA_signal_16989 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16993 ;
    wire new_AGEMA_signal_16994 ;
    wire new_AGEMA_signal_16995 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_16999 ;
    wire new_AGEMA_signal_17000 ;
    wire new_AGEMA_signal_17001 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire new_AGEMA_signal_17005 ;
    wire new_AGEMA_signal_17006 ;
    wire new_AGEMA_signal_17007 ;
    wire new_AGEMA_signal_17008 ;
    wire new_AGEMA_signal_17009 ;
    wire new_AGEMA_signal_17010 ;
    wire new_AGEMA_signal_17011 ;
    wire new_AGEMA_signal_17012 ;
    wire new_AGEMA_signal_17013 ;
    wire new_AGEMA_signal_17014 ;
    wire new_AGEMA_signal_17015 ;
    wire new_AGEMA_signal_17016 ;
    wire new_AGEMA_signal_17017 ;
    wire new_AGEMA_signal_17018 ;
    wire new_AGEMA_signal_17019 ;
    wire new_AGEMA_signal_17020 ;
    wire new_AGEMA_signal_17021 ;
    wire new_AGEMA_signal_17022 ;
    wire new_AGEMA_signal_17023 ;
    wire new_AGEMA_signal_17024 ;
    wire new_AGEMA_signal_17025 ;
    wire new_AGEMA_signal_17026 ;
    wire new_AGEMA_signal_17027 ;
    wire new_AGEMA_signal_17028 ;
    wire new_AGEMA_signal_17029 ;
    wire new_AGEMA_signal_17030 ;
    wire new_AGEMA_signal_17031 ;
    wire new_AGEMA_signal_17032 ;
    wire new_AGEMA_signal_17033 ;
    wire new_AGEMA_signal_17034 ;
    wire new_AGEMA_signal_17035 ;
    wire new_AGEMA_signal_17036 ;
    wire new_AGEMA_signal_17037 ;
    wire new_AGEMA_signal_17038 ;
    wire new_AGEMA_signal_17039 ;
    wire new_AGEMA_signal_17040 ;
    wire new_AGEMA_signal_17041 ;
    wire new_AGEMA_signal_17042 ;
    wire new_AGEMA_signal_17043 ;
    wire new_AGEMA_signal_17044 ;
    wire new_AGEMA_signal_17045 ;
    wire new_AGEMA_signal_17046 ;
    wire new_AGEMA_signal_17047 ;
    wire new_AGEMA_signal_17048 ;
    wire new_AGEMA_signal_17049 ;
    wire new_AGEMA_signal_17050 ;
    wire new_AGEMA_signal_17051 ;
    wire new_AGEMA_signal_17052 ;
    wire new_AGEMA_signal_17053 ;
    wire new_AGEMA_signal_17054 ;
    wire new_AGEMA_signal_17055 ;
    wire new_AGEMA_signal_17056 ;
    wire new_AGEMA_signal_17057 ;
    wire new_AGEMA_signal_17058 ;
    wire new_AGEMA_signal_17059 ;
    wire new_AGEMA_signal_17060 ;
    wire new_AGEMA_signal_17061 ;
    wire new_AGEMA_signal_17062 ;
    wire new_AGEMA_signal_17063 ;
    wire new_AGEMA_signal_17064 ;
    wire new_AGEMA_signal_17065 ;
    wire new_AGEMA_signal_17066 ;
    wire new_AGEMA_signal_17067 ;
    wire new_AGEMA_signal_17068 ;
    wire new_AGEMA_signal_17069 ;
    wire new_AGEMA_signal_17070 ;
    wire new_AGEMA_signal_17071 ;
    wire new_AGEMA_signal_17072 ;
    wire new_AGEMA_signal_17073 ;
    wire new_AGEMA_signal_17074 ;
    wire new_AGEMA_signal_17075 ;
    wire new_AGEMA_signal_17076 ;
    wire new_AGEMA_signal_17077 ;
    wire new_AGEMA_signal_17078 ;
    wire new_AGEMA_signal_17079 ;
    wire new_AGEMA_signal_17080 ;
    wire new_AGEMA_signal_17081 ;
    wire new_AGEMA_signal_17082 ;
    wire new_AGEMA_signal_17083 ;
    wire new_AGEMA_signal_17084 ;
    wire new_AGEMA_signal_17085 ;
    wire new_AGEMA_signal_17086 ;
    wire new_AGEMA_signal_17087 ;
    wire new_AGEMA_signal_17088 ;
    wire new_AGEMA_signal_17089 ;
    wire new_AGEMA_signal_17090 ;
    wire new_AGEMA_signal_17091 ;
    wire new_AGEMA_signal_17092 ;
    wire new_AGEMA_signal_17093 ;
    wire new_AGEMA_signal_17094 ;
    wire new_AGEMA_signal_17095 ;
    wire new_AGEMA_signal_17096 ;
    wire new_AGEMA_signal_17097 ;
    wire new_AGEMA_signal_17098 ;
    wire new_AGEMA_signal_17099 ;
    wire new_AGEMA_signal_17100 ;
    wire new_AGEMA_signal_17101 ;
    wire new_AGEMA_signal_17102 ;
    wire new_AGEMA_signal_17103 ;
    wire new_AGEMA_signal_17104 ;
    wire new_AGEMA_signal_17105 ;
    wire new_AGEMA_signal_17106 ;
    wire new_AGEMA_signal_17107 ;
    wire new_AGEMA_signal_17108 ;
    wire new_AGEMA_signal_17109 ;
    wire new_AGEMA_signal_17110 ;
    wire new_AGEMA_signal_17111 ;
    wire new_AGEMA_signal_17112 ;
    wire new_AGEMA_signal_17113 ;
    wire new_AGEMA_signal_17114 ;
    wire new_AGEMA_signal_17115 ;
    wire new_AGEMA_signal_17116 ;
    wire new_AGEMA_signal_17117 ;
    wire new_AGEMA_signal_17118 ;
    wire new_AGEMA_signal_17119 ;
    wire new_AGEMA_signal_17120 ;
    wire new_AGEMA_signal_17121 ;
    wire new_AGEMA_signal_17122 ;
    wire new_AGEMA_signal_17123 ;
    wire new_AGEMA_signal_17124 ;
    wire new_AGEMA_signal_17125 ;
    wire new_AGEMA_signal_17126 ;
    wire new_AGEMA_signal_17127 ;
    wire new_AGEMA_signal_17128 ;
    wire new_AGEMA_signal_17129 ;
    wire new_AGEMA_signal_17130 ;
    wire new_AGEMA_signal_17131 ;
    wire new_AGEMA_signal_17132 ;
    wire new_AGEMA_signal_17133 ;
    wire new_AGEMA_signal_17134 ;
    wire new_AGEMA_signal_17135 ;
    wire new_AGEMA_signal_17136 ;
    wire new_AGEMA_signal_17137 ;
    wire new_AGEMA_signal_17138 ;
    wire new_AGEMA_signal_17139 ;
    wire new_AGEMA_signal_17140 ;
    wire new_AGEMA_signal_17141 ;
    wire new_AGEMA_signal_17142 ;
    wire new_AGEMA_signal_17143 ;
    wire new_AGEMA_signal_17144 ;
    wire new_AGEMA_signal_17145 ;
    wire new_AGEMA_signal_17146 ;
    wire new_AGEMA_signal_17147 ;
    wire new_AGEMA_signal_17148 ;
    wire new_AGEMA_signal_17149 ;
    wire new_AGEMA_signal_17150 ;
    wire new_AGEMA_signal_17151 ;
    wire new_AGEMA_signal_17152 ;
    wire new_AGEMA_signal_17153 ;
    wire new_AGEMA_signal_17154 ;
    wire new_AGEMA_signal_17155 ;
    wire new_AGEMA_signal_17156 ;
    wire new_AGEMA_signal_17157 ;
    wire new_AGEMA_signal_17158 ;
    wire new_AGEMA_signal_17159 ;
    wire new_AGEMA_signal_17160 ;
    wire new_AGEMA_signal_17161 ;
    wire new_AGEMA_signal_17162 ;
    wire new_AGEMA_signal_17163 ;
    wire new_AGEMA_signal_17164 ;
    wire new_AGEMA_signal_17165 ;
    wire new_AGEMA_signal_17166 ;
    wire new_AGEMA_signal_17167 ;
    wire new_AGEMA_signal_17168 ;
    wire new_AGEMA_signal_17169 ;
    wire new_AGEMA_signal_17170 ;
    wire new_AGEMA_signal_17171 ;
    wire new_AGEMA_signal_17172 ;
    wire new_AGEMA_signal_17173 ;
    wire new_AGEMA_signal_17174 ;
    wire new_AGEMA_signal_17175 ;
    wire new_AGEMA_signal_17176 ;
    wire new_AGEMA_signal_17177 ;
    wire new_AGEMA_signal_17178 ;
    wire new_AGEMA_signal_17179 ;
    wire new_AGEMA_signal_17180 ;
    wire new_AGEMA_signal_17181 ;
    wire new_AGEMA_signal_17182 ;
    wire new_AGEMA_signal_17183 ;
    wire new_AGEMA_signal_17184 ;
    wire new_AGEMA_signal_17185 ;
    wire new_AGEMA_signal_17186 ;
    wire new_AGEMA_signal_17187 ;
    wire new_AGEMA_signal_17188 ;
    wire new_AGEMA_signal_17189 ;
    wire new_AGEMA_signal_17190 ;
    wire new_AGEMA_signal_17191 ;
    wire new_AGEMA_signal_17192 ;
    wire new_AGEMA_signal_17193 ;
    wire new_AGEMA_signal_17194 ;
    wire new_AGEMA_signal_17195 ;
    wire new_AGEMA_signal_17196 ;
    wire new_AGEMA_signal_17197 ;
    wire new_AGEMA_signal_17198 ;
    wire new_AGEMA_signal_17199 ;
    wire new_AGEMA_signal_17200 ;
    wire new_AGEMA_signal_17201 ;
    wire new_AGEMA_signal_17202 ;
    wire new_AGEMA_signal_17203 ;
    wire new_AGEMA_signal_17204 ;
    wire new_AGEMA_signal_17205 ;
    wire new_AGEMA_signal_17206 ;
    wire new_AGEMA_signal_17207 ;
    wire new_AGEMA_signal_17208 ;
    wire new_AGEMA_signal_17209 ;
    wire new_AGEMA_signal_17210 ;
    wire new_AGEMA_signal_17211 ;
    wire new_AGEMA_signal_17212 ;
    wire new_AGEMA_signal_17213 ;
    wire new_AGEMA_signal_17214 ;
    wire new_AGEMA_signal_17215 ;
    wire new_AGEMA_signal_17216 ;
    wire new_AGEMA_signal_17217 ;
    wire new_AGEMA_signal_17218 ;
    wire new_AGEMA_signal_17219 ;
    wire new_AGEMA_signal_17220 ;
    wire new_AGEMA_signal_17221 ;
    wire new_AGEMA_signal_17222 ;
    wire new_AGEMA_signal_17223 ;
    wire new_AGEMA_signal_17224 ;
    wire new_AGEMA_signal_17225 ;
    wire new_AGEMA_signal_17226 ;
    wire new_AGEMA_signal_17227 ;
    wire new_AGEMA_signal_17228 ;
    wire new_AGEMA_signal_17229 ;
    wire new_AGEMA_signal_17230 ;
    wire new_AGEMA_signal_17231 ;
    wire new_AGEMA_signal_17232 ;
    wire new_AGEMA_signal_17233 ;
    wire new_AGEMA_signal_17234 ;
    wire new_AGEMA_signal_17235 ;
    wire new_AGEMA_signal_17236 ;
    wire new_AGEMA_signal_17237 ;
    wire new_AGEMA_signal_17238 ;
    wire new_AGEMA_signal_17239 ;
    wire new_AGEMA_signal_17240 ;
    wire new_AGEMA_signal_17241 ;
    wire new_AGEMA_signal_17242 ;
    wire new_AGEMA_signal_17243 ;
    wire new_AGEMA_signal_17244 ;
    wire new_AGEMA_signal_17245 ;
    wire new_AGEMA_signal_17246 ;
    wire new_AGEMA_signal_17247 ;
    wire new_AGEMA_signal_17248 ;
    wire new_AGEMA_signal_17249 ;
    wire new_AGEMA_signal_17250 ;
    wire new_AGEMA_signal_17251 ;
    wire new_AGEMA_signal_17252 ;
    wire new_AGEMA_signal_17253 ;
    wire new_AGEMA_signal_17254 ;
    wire new_AGEMA_signal_17255 ;
    wire new_AGEMA_signal_17256 ;
    wire new_AGEMA_signal_17257 ;
    wire new_AGEMA_signal_17258 ;
    wire new_AGEMA_signal_17259 ;
    wire new_AGEMA_signal_17260 ;
    wire new_AGEMA_signal_17261 ;
    wire new_AGEMA_signal_17262 ;
    wire new_AGEMA_signal_17263 ;
    wire new_AGEMA_signal_17264 ;
    wire new_AGEMA_signal_17265 ;
    wire new_AGEMA_signal_17266 ;
    wire new_AGEMA_signal_17267 ;
    wire new_AGEMA_signal_17268 ;
    wire new_AGEMA_signal_17269 ;
    wire new_AGEMA_signal_17270 ;
    wire new_AGEMA_signal_17271 ;
    wire new_AGEMA_signal_17272 ;
    wire new_AGEMA_signal_17273 ;
    wire new_AGEMA_signal_17274 ;
    wire new_AGEMA_signal_17275 ;
    wire new_AGEMA_signal_17276 ;
    wire new_AGEMA_signal_17277 ;
    wire new_AGEMA_signal_17278 ;
    wire new_AGEMA_signal_17279 ;
    wire new_AGEMA_signal_17280 ;
    wire new_AGEMA_signal_17281 ;
    wire new_AGEMA_signal_17282 ;
    wire new_AGEMA_signal_17283 ;
    wire new_AGEMA_signal_17284 ;
    wire new_AGEMA_signal_17285 ;
    wire new_AGEMA_signal_17286 ;
    wire new_AGEMA_signal_17287 ;
    wire new_AGEMA_signal_17288 ;
    wire new_AGEMA_signal_17289 ;
    wire new_AGEMA_signal_17290 ;
    wire new_AGEMA_signal_17291 ;
    wire new_AGEMA_signal_17292 ;
    wire new_AGEMA_signal_17293 ;
    wire new_AGEMA_signal_17294 ;
    wire new_AGEMA_signal_17295 ;
    wire new_AGEMA_signal_17296 ;
    wire new_AGEMA_signal_17297 ;
    wire new_AGEMA_signal_17298 ;
    wire new_AGEMA_signal_17299 ;
    wire new_AGEMA_signal_17300 ;
    wire new_AGEMA_signal_17301 ;
    wire new_AGEMA_signal_17302 ;
    wire new_AGEMA_signal_17303 ;
    wire new_AGEMA_signal_17304 ;
    wire new_AGEMA_signal_17305 ;
    wire new_AGEMA_signal_17306 ;
    wire new_AGEMA_signal_17307 ;
    wire new_AGEMA_signal_17308 ;
    wire new_AGEMA_signal_17309 ;
    wire new_AGEMA_signal_17310 ;
    wire new_AGEMA_signal_17311 ;
    wire new_AGEMA_signal_17312 ;
    wire new_AGEMA_signal_17313 ;
    wire new_AGEMA_signal_17314 ;
    wire new_AGEMA_signal_17315 ;
    wire new_AGEMA_signal_17316 ;
    wire new_AGEMA_signal_17317 ;
    wire new_AGEMA_signal_17318 ;
    wire new_AGEMA_signal_17319 ;
    wire new_AGEMA_signal_17320 ;
    wire new_AGEMA_signal_17321 ;
    wire new_AGEMA_signal_17322 ;
    wire new_AGEMA_signal_17323 ;
    wire new_AGEMA_signal_17324 ;
    wire new_AGEMA_signal_17325 ;
    wire new_AGEMA_signal_17326 ;
    wire new_AGEMA_signal_17327 ;
    wire new_AGEMA_signal_17328 ;
    wire new_AGEMA_signal_17329 ;
    wire new_AGEMA_signal_17330 ;
    wire new_AGEMA_signal_17331 ;
    wire new_AGEMA_signal_17332 ;
    wire new_AGEMA_signal_17333 ;
    wire new_AGEMA_signal_17334 ;
    wire new_AGEMA_signal_17335 ;
    wire new_AGEMA_signal_17336 ;
    wire new_AGEMA_signal_17337 ;
    wire new_AGEMA_signal_17338 ;
    wire new_AGEMA_signal_17339 ;
    wire new_AGEMA_signal_17340 ;
    wire new_AGEMA_signal_17341 ;
    wire new_AGEMA_signal_17342 ;
    wire new_AGEMA_signal_17343 ;
    wire new_AGEMA_signal_17344 ;
    wire new_AGEMA_signal_17345 ;
    wire new_AGEMA_signal_17346 ;
    wire new_AGEMA_signal_17347 ;
    wire new_AGEMA_signal_17348 ;
    wire new_AGEMA_signal_17349 ;
    wire new_AGEMA_signal_17350 ;
    wire new_AGEMA_signal_17351 ;
    wire new_AGEMA_signal_17352 ;
    wire new_AGEMA_signal_17353 ;
    wire new_AGEMA_signal_17354 ;
    wire new_AGEMA_signal_17355 ;
    wire new_AGEMA_signal_17356 ;
    wire new_AGEMA_signal_17357 ;
    wire new_AGEMA_signal_17358 ;
    wire new_AGEMA_signal_17359 ;
    wire new_AGEMA_signal_17360 ;
    wire new_AGEMA_signal_17361 ;
    wire new_AGEMA_signal_17362 ;
    wire new_AGEMA_signal_17363 ;
    wire new_AGEMA_signal_17364 ;
    wire new_AGEMA_signal_17365 ;
    wire new_AGEMA_signal_17366 ;
    wire new_AGEMA_signal_17367 ;
    wire new_AGEMA_signal_17368 ;
    wire new_AGEMA_signal_17369 ;
    wire new_AGEMA_signal_17370 ;
    wire new_AGEMA_signal_17371 ;
    wire new_AGEMA_signal_17372 ;
    wire new_AGEMA_signal_17373 ;
    wire new_AGEMA_signal_17374 ;
    wire new_AGEMA_signal_17375 ;
    wire new_AGEMA_signal_17376 ;
    wire new_AGEMA_signal_17377 ;
    wire new_AGEMA_signal_17378 ;
    wire new_AGEMA_signal_17379 ;
    wire new_AGEMA_signal_17380 ;
    wire new_AGEMA_signal_17381 ;
    wire new_AGEMA_signal_17382 ;
    wire new_AGEMA_signal_17383 ;
    wire new_AGEMA_signal_17384 ;
    wire new_AGEMA_signal_17385 ;
    wire new_AGEMA_signal_17386 ;
    wire new_AGEMA_signal_17387 ;
    wire new_AGEMA_signal_17388 ;
    wire new_AGEMA_signal_17389 ;
    wire new_AGEMA_signal_17390 ;
    wire new_AGEMA_signal_17391 ;
    wire new_AGEMA_signal_17392 ;
    wire new_AGEMA_signal_17393 ;
    wire new_AGEMA_signal_17394 ;
    wire new_AGEMA_signal_17395 ;
    wire new_AGEMA_signal_17396 ;
    wire new_AGEMA_signal_17397 ;
    wire new_AGEMA_signal_17398 ;
    wire new_AGEMA_signal_17399 ;
    wire new_AGEMA_signal_17400 ;
    wire new_AGEMA_signal_17401 ;
    wire new_AGEMA_signal_17402 ;
    wire new_AGEMA_signal_17403 ;
    wire new_AGEMA_signal_17404 ;
    wire new_AGEMA_signal_17405 ;
    wire new_AGEMA_signal_17406 ;
    wire new_AGEMA_signal_17407 ;
    wire new_AGEMA_signal_17408 ;
    wire new_AGEMA_signal_17409 ;
    wire new_AGEMA_signal_17410 ;
    wire new_AGEMA_signal_17411 ;
    wire new_AGEMA_signal_17412 ;
    wire new_AGEMA_signal_17413 ;
    wire new_AGEMA_signal_17414 ;
    wire new_AGEMA_signal_17415 ;
    wire new_AGEMA_signal_17416 ;
    wire new_AGEMA_signal_17417 ;
    wire new_AGEMA_signal_17418 ;
    wire new_AGEMA_signal_17419 ;
    wire new_AGEMA_signal_17420 ;
    wire new_AGEMA_signal_17421 ;
    wire new_AGEMA_signal_17422 ;
    wire new_AGEMA_signal_17423 ;
    wire new_AGEMA_signal_17424 ;
    wire new_AGEMA_signal_17425 ;
    wire new_AGEMA_signal_17426 ;
    wire new_AGEMA_signal_17427 ;
    wire new_AGEMA_signal_17428 ;
    wire new_AGEMA_signal_17429 ;
    wire new_AGEMA_signal_17430 ;
    wire new_AGEMA_signal_17431 ;
    wire new_AGEMA_signal_17432 ;
    wire new_AGEMA_signal_17433 ;
    wire new_AGEMA_signal_17434 ;
    wire new_AGEMA_signal_17435 ;
    wire new_AGEMA_signal_17436 ;
    wire new_AGEMA_signal_17437 ;
    wire new_AGEMA_signal_17438 ;
    wire new_AGEMA_signal_17439 ;
    wire new_AGEMA_signal_17440 ;
    wire new_AGEMA_signal_17441 ;
    wire new_AGEMA_signal_17442 ;
    wire new_AGEMA_signal_17443 ;
    wire new_AGEMA_signal_17444 ;
    wire new_AGEMA_signal_17445 ;
    wire new_AGEMA_signal_17446 ;
    wire new_AGEMA_signal_17447 ;
    wire new_AGEMA_signal_17448 ;
    wire new_AGEMA_signal_17449 ;
    wire new_AGEMA_signal_17450 ;
    wire new_AGEMA_signal_17451 ;
    wire new_AGEMA_signal_17452 ;
    wire new_AGEMA_signal_17453 ;
    wire new_AGEMA_signal_17454 ;
    wire new_AGEMA_signal_17455 ;
    wire new_AGEMA_signal_17456 ;
    wire new_AGEMA_signal_17457 ;
    wire new_AGEMA_signal_17458 ;
    wire new_AGEMA_signal_17459 ;
    wire new_AGEMA_signal_17460 ;
    wire new_AGEMA_signal_17461 ;
    wire new_AGEMA_signal_17462 ;
    wire new_AGEMA_signal_17463 ;
    wire new_AGEMA_signal_17464 ;
    wire new_AGEMA_signal_17465 ;
    wire new_AGEMA_signal_17466 ;
    wire new_AGEMA_signal_17467 ;
    wire new_AGEMA_signal_17468 ;
    wire new_AGEMA_signal_17469 ;
    wire new_AGEMA_signal_17470 ;
    wire new_AGEMA_signal_17471 ;
    wire new_AGEMA_signal_17472 ;
    wire new_AGEMA_signal_17473 ;
    wire new_AGEMA_signal_17474 ;
    wire new_AGEMA_signal_17475 ;
    wire new_AGEMA_signal_17476 ;
    wire new_AGEMA_signal_17477 ;
    wire new_AGEMA_signal_17478 ;
    wire new_AGEMA_signal_17479 ;
    wire new_AGEMA_signal_17480 ;
    wire new_AGEMA_signal_17481 ;
    wire new_AGEMA_signal_17482 ;
    wire new_AGEMA_signal_17483 ;
    wire new_AGEMA_signal_17484 ;
    wire new_AGEMA_signal_17485 ;
    wire new_AGEMA_signal_17486 ;
    wire new_AGEMA_signal_17487 ;
    wire new_AGEMA_signal_17488 ;
    wire new_AGEMA_signal_17489 ;
    wire new_AGEMA_signal_17490 ;
    wire new_AGEMA_signal_17491 ;
    wire new_AGEMA_signal_17492 ;
    wire new_AGEMA_signal_17493 ;
    wire new_AGEMA_signal_17494 ;
    wire new_AGEMA_signal_17495 ;
    wire new_AGEMA_signal_17496 ;
    wire new_AGEMA_signal_17497 ;
    wire new_AGEMA_signal_17498 ;
    wire new_AGEMA_signal_17499 ;
    wire new_AGEMA_signal_17500 ;
    wire new_AGEMA_signal_17501 ;
    wire new_AGEMA_signal_17502 ;
    wire new_AGEMA_signal_17503 ;
    wire new_AGEMA_signal_17504 ;
    wire new_AGEMA_signal_17505 ;
    wire new_AGEMA_signal_17506 ;
    wire new_AGEMA_signal_17507 ;
    wire new_AGEMA_signal_17508 ;
    wire new_AGEMA_signal_17509 ;
    wire new_AGEMA_signal_17510 ;
    wire new_AGEMA_signal_17511 ;
    wire new_AGEMA_signal_17512 ;
    wire new_AGEMA_signal_17513 ;
    wire new_AGEMA_signal_17514 ;
    wire new_AGEMA_signal_17515 ;
    wire new_AGEMA_signal_17516 ;
    wire new_AGEMA_signal_17517 ;
    wire new_AGEMA_signal_17518 ;
    wire new_AGEMA_signal_17519 ;
    wire new_AGEMA_signal_17520 ;
    wire new_AGEMA_signal_17521 ;
    wire new_AGEMA_signal_17522 ;
    wire new_AGEMA_signal_17523 ;
    wire new_AGEMA_signal_17524 ;
    wire new_AGEMA_signal_17525 ;
    wire new_AGEMA_signal_17526 ;
    wire new_AGEMA_signal_17527 ;
    wire new_AGEMA_signal_17528 ;
    wire new_AGEMA_signal_17529 ;
    wire new_AGEMA_signal_17530 ;
    wire new_AGEMA_signal_17531 ;
    wire new_AGEMA_signal_17532 ;
    wire new_AGEMA_signal_17533 ;
    wire new_AGEMA_signal_17534 ;
    wire new_AGEMA_signal_17535 ;
    wire new_AGEMA_signal_17536 ;
    wire new_AGEMA_signal_17537 ;
    wire new_AGEMA_signal_17538 ;
    wire new_AGEMA_signal_17539 ;
    wire new_AGEMA_signal_17540 ;
    wire new_AGEMA_signal_17541 ;
    wire new_AGEMA_signal_17542 ;
    wire new_AGEMA_signal_17543 ;
    wire new_AGEMA_signal_17544 ;
    wire new_AGEMA_signal_17545 ;
    wire new_AGEMA_signal_17546 ;
    wire new_AGEMA_signal_17547 ;
    wire new_AGEMA_signal_17548 ;
    wire new_AGEMA_signal_17549 ;
    wire new_AGEMA_signal_17550 ;
    wire new_AGEMA_signal_17551 ;
    wire new_AGEMA_signal_17552 ;
    wire new_AGEMA_signal_17553 ;
    wire new_AGEMA_signal_17554 ;
    wire new_AGEMA_signal_17555 ;
    wire new_AGEMA_signal_17556 ;
    wire new_AGEMA_signal_17557 ;
    wire new_AGEMA_signal_17558 ;
    wire new_AGEMA_signal_17559 ;
    wire new_AGEMA_signal_17560 ;
    wire new_AGEMA_signal_17561 ;
    wire new_AGEMA_signal_17562 ;
    wire new_AGEMA_signal_17563 ;
    wire new_AGEMA_signal_17564 ;
    wire new_AGEMA_signal_17565 ;
    wire new_AGEMA_signal_17566 ;
    wire new_AGEMA_signal_17567 ;
    wire new_AGEMA_signal_17568 ;
    wire new_AGEMA_signal_17569 ;
    wire new_AGEMA_signal_17570 ;
    wire new_AGEMA_signal_17571 ;
    wire new_AGEMA_signal_17572 ;
    wire new_AGEMA_signal_17573 ;
    wire new_AGEMA_signal_17574 ;
    wire new_AGEMA_signal_17575 ;
    wire new_AGEMA_signal_17576 ;
    wire new_AGEMA_signal_17577 ;
    wire new_AGEMA_signal_17578 ;
    wire new_AGEMA_signal_17579 ;
    wire new_AGEMA_signal_17580 ;
    wire new_AGEMA_signal_17581 ;
    wire new_AGEMA_signal_17582 ;
    wire new_AGEMA_signal_17583 ;
    wire new_AGEMA_signal_17584 ;
    wire new_AGEMA_signal_17585 ;
    wire new_AGEMA_signal_17586 ;
    wire new_AGEMA_signal_17587 ;
    wire new_AGEMA_signal_17588 ;
    wire new_AGEMA_signal_17589 ;
    wire new_AGEMA_signal_17590 ;
    wire new_AGEMA_signal_17591 ;
    wire new_AGEMA_signal_17592 ;
    wire new_AGEMA_signal_17593 ;
    wire new_AGEMA_signal_17594 ;
    wire new_AGEMA_signal_17595 ;
    wire new_AGEMA_signal_17596 ;
    wire new_AGEMA_signal_17597 ;
    wire new_AGEMA_signal_17598 ;
    wire new_AGEMA_signal_17599 ;
    wire new_AGEMA_signal_17600 ;
    wire new_AGEMA_signal_17601 ;
    wire new_AGEMA_signal_17602 ;
    wire new_AGEMA_signal_17603 ;
    wire new_AGEMA_signal_17604 ;
    wire new_AGEMA_signal_17605 ;
    wire new_AGEMA_signal_17606 ;
    wire new_AGEMA_signal_17607 ;
    wire new_AGEMA_signal_17608 ;
    wire new_AGEMA_signal_17609 ;
    wire new_AGEMA_signal_17610 ;
    wire new_AGEMA_signal_17611 ;
    wire new_AGEMA_signal_17612 ;
    wire new_AGEMA_signal_17613 ;
    wire new_AGEMA_signal_17614 ;
    wire new_AGEMA_signal_17615 ;
    wire new_AGEMA_signal_17616 ;
    wire new_AGEMA_signal_17617 ;
    wire new_AGEMA_signal_17618 ;
    wire new_AGEMA_signal_17619 ;
    wire new_AGEMA_signal_17620 ;
    wire new_AGEMA_signal_17621 ;
    wire new_AGEMA_signal_17622 ;
    wire new_AGEMA_signal_17623 ;
    wire new_AGEMA_signal_17624 ;
    wire new_AGEMA_signal_17625 ;
    wire new_AGEMA_signal_17626 ;
    wire new_AGEMA_signal_17627 ;
    wire new_AGEMA_signal_17628 ;
    wire new_AGEMA_signal_17629 ;
    wire new_AGEMA_signal_17630 ;
    wire new_AGEMA_signal_17631 ;
    wire new_AGEMA_signal_17632 ;
    wire new_AGEMA_signal_17633 ;
    wire new_AGEMA_signal_17634 ;
    wire new_AGEMA_signal_17635 ;
    wire new_AGEMA_signal_17636 ;
    wire new_AGEMA_signal_17637 ;
    wire new_AGEMA_signal_17638 ;
    wire new_AGEMA_signal_17639 ;
    wire new_AGEMA_signal_17640 ;
    wire new_AGEMA_signal_17641 ;
    wire new_AGEMA_signal_17642 ;
    wire new_AGEMA_signal_17643 ;
    wire new_AGEMA_signal_17644 ;
    wire new_AGEMA_signal_17645 ;
    wire new_AGEMA_signal_17646 ;
    wire new_AGEMA_signal_17647 ;
    wire new_AGEMA_signal_17648 ;
    wire new_AGEMA_signal_17649 ;
    wire new_AGEMA_signal_17650 ;
    wire new_AGEMA_signal_17651 ;
    wire new_AGEMA_signal_17652 ;
    wire new_AGEMA_signal_17653 ;
    wire new_AGEMA_signal_17654 ;
    wire new_AGEMA_signal_17655 ;
    wire new_AGEMA_signal_17656 ;
    wire new_AGEMA_signal_17657 ;
    wire new_AGEMA_signal_17658 ;
    wire new_AGEMA_signal_17659 ;
    wire new_AGEMA_signal_17660 ;
    wire new_AGEMA_signal_17661 ;
    wire new_AGEMA_signal_17662 ;
    wire new_AGEMA_signal_17663 ;
    wire new_AGEMA_signal_17664 ;
    wire new_AGEMA_signal_17665 ;
    wire new_AGEMA_signal_17666 ;
    wire new_AGEMA_signal_17667 ;
    wire new_AGEMA_signal_17668 ;
    wire new_AGEMA_signal_17669 ;
    wire new_AGEMA_signal_17670 ;
    wire new_AGEMA_signal_17671 ;
    wire new_AGEMA_signal_17672 ;
    wire new_AGEMA_signal_17673 ;
    wire new_AGEMA_signal_17674 ;
    wire new_AGEMA_signal_17675 ;
    wire new_AGEMA_signal_17676 ;
    wire new_AGEMA_signal_17677 ;
    wire new_AGEMA_signal_17678 ;
    wire new_AGEMA_signal_17679 ;
    wire new_AGEMA_signal_17680 ;
    wire new_AGEMA_signal_17681 ;
    wire new_AGEMA_signal_17682 ;
    wire new_AGEMA_signal_17683 ;
    wire new_AGEMA_signal_17684 ;
    wire new_AGEMA_signal_17685 ;
    wire new_AGEMA_signal_17686 ;
    wire new_AGEMA_signal_17687 ;
    wire new_AGEMA_signal_17688 ;
    wire new_AGEMA_signal_17689 ;
    wire new_AGEMA_signal_17690 ;
    wire new_AGEMA_signal_17691 ;
    wire new_AGEMA_signal_17692 ;
    wire new_AGEMA_signal_17693 ;
    wire new_AGEMA_signal_17694 ;
    wire new_AGEMA_signal_17695 ;
    wire new_AGEMA_signal_17696 ;
    wire new_AGEMA_signal_17697 ;
    wire new_AGEMA_signal_17698 ;
    wire new_AGEMA_signal_17699 ;
    wire new_AGEMA_signal_17700 ;
    wire new_AGEMA_signal_17701 ;
    wire new_AGEMA_signal_17702 ;
    wire new_AGEMA_signal_17703 ;
    wire new_AGEMA_signal_17704 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17708 ;
    wire new_AGEMA_signal_17709 ;
    wire new_AGEMA_signal_17710 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17714 ;
    wire new_AGEMA_signal_17715 ;
    wire new_AGEMA_signal_17716 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17720 ;
    wire new_AGEMA_signal_17721 ;
    wire new_AGEMA_signal_17722 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17726 ;
    wire new_AGEMA_signal_17727 ;
    wire new_AGEMA_signal_17728 ;
    wire new_AGEMA_signal_17729 ;
    wire new_AGEMA_signal_17730 ;
    wire new_AGEMA_signal_17731 ;
    wire new_AGEMA_signal_17732 ;
    wire new_AGEMA_signal_17733 ;
    wire new_AGEMA_signal_17734 ;
    wire new_AGEMA_signal_17735 ;
    wire new_AGEMA_signal_17736 ;
    wire new_AGEMA_signal_17737 ;
    wire new_AGEMA_signal_17738 ;
    wire new_AGEMA_signal_17739 ;
    wire new_AGEMA_signal_17740 ;
    wire new_AGEMA_signal_17741 ;
    wire new_AGEMA_signal_17742 ;
    wire new_AGEMA_signal_17743 ;
    wire new_AGEMA_signal_17744 ;
    wire new_AGEMA_signal_17745 ;
    wire new_AGEMA_signal_17746 ;
    wire new_AGEMA_signal_17747 ;
    wire new_AGEMA_signal_17748 ;
    wire new_AGEMA_signal_17749 ;
    wire new_AGEMA_signal_17750 ;
    wire new_AGEMA_signal_17751 ;
    wire new_AGEMA_signal_17752 ;
    wire new_AGEMA_signal_17753 ;
    wire new_AGEMA_signal_17754 ;
    wire new_AGEMA_signal_17755 ;
    wire new_AGEMA_signal_17756 ;
    wire new_AGEMA_signal_17757 ;
    wire new_AGEMA_signal_17758 ;
    wire new_AGEMA_signal_17759 ;
    wire new_AGEMA_signal_17760 ;
    wire new_AGEMA_signal_17761 ;
    wire new_AGEMA_signal_17762 ;
    wire new_AGEMA_signal_17763 ;
    wire new_AGEMA_signal_17764 ;
    wire new_AGEMA_signal_17765 ;
    wire new_AGEMA_signal_17766 ;
    wire new_AGEMA_signal_17767 ;
    wire new_AGEMA_signal_17768 ;
    wire new_AGEMA_signal_17769 ;
    wire new_AGEMA_signal_17770 ;
    wire new_AGEMA_signal_17771 ;
    wire new_AGEMA_signal_17772 ;
    wire new_AGEMA_signal_17773 ;
    wire new_AGEMA_signal_17774 ;
    wire new_AGEMA_signal_17775 ;
    wire new_AGEMA_signal_17776 ;
    wire new_AGEMA_signal_17777 ;
    wire new_AGEMA_signal_17778 ;
    wire new_AGEMA_signal_17779 ;
    wire new_AGEMA_signal_17780 ;
    wire new_AGEMA_signal_17781 ;
    wire new_AGEMA_signal_17782 ;
    wire new_AGEMA_signal_17783 ;
    wire new_AGEMA_signal_17784 ;
    wire new_AGEMA_signal_17785 ;
    wire new_AGEMA_signal_17786 ;
    wire new_AGEMA_signal_17787 ;
    wire new_AGEMA_signal_17788 ;
    wire new_AGEMA_signal_17789 ;
    wire new_AGEMA_signal_17790 ;
    wire new_AGEMA_signal_17791 ;
    wire new_AGEMA_signal_17792 ;
    wire new_AGEMA_signal_17793 ;
    wire new_AGEMA_signal_17794 ;
    wire new_AGEMA_signal_17795 ;
    wire new_AGEMA_signal_17796 ;
    wire new_AGEMA_signal_17797 ;
    wire new_AGEMA_signal_17798 ;
    wire new_AGEMA_signal_17799 ;
    wire new_AGEMA_signal_17800 ;
    wire new_AGEMA_signal_17801 ;
    wire new_AGEMA_signal_17802 ;
    wire new_AGEMA_signal_17803 ;
    wire new_AGEMA_signal_17804 ;
    wire new_AGEMA_signal_17805 ;
    wire new_AGEMA_signal_17806 ;
    wire new_AGEMA_signal_17807 ;
    wire new_AGEMA_signal_17808 ;
    wire new_AGEMA_signal_17809 ;
    wire new_AGEMA_signal_17810 ;
    wire new_AGEMA_signal_17811 ;
    wire new_AGEMA_signal_17812 ;
    wire new_AGEMA_signal_17813 ;
    wire new_AGEMA_signal_17814 ;
    wire new_AGEMA_signal_17815 ;
    wire new_AGEMA_signal_17816 ;
    wire new_AGEMA_signal_17817 ;
    wire new_AGEMA_signal_17818 ;
    wire new_AGEMA_signal_17819 ;
    wire new_AGEMA_signal_17820 ;
    wire new_AGEMA_signal_17821 ;
    wire new_AGEMA_signal_17822 ;
    wire new_AGEMA_signal_17823 ;
    wire new_AGEMA_signal_17824 ;
    wire new_AGEMA_signal_17825 ;
    wire new_AGEMA_signal_17826 ;
    wire new_AGEMA_signal_17827 ;
    wire new_AGEMA_signal_17828 ;
    wire new_AGEMA_signal_17829 ;
    wire new_AGEMA_signal_17830 ;
    wire new_AGEMA_signal_17831 ;
    wire new_AGEMA_signal_17832 ;
    wire new_AGEMA_signal_17833 ;
    wire new_AGEMA_signal_17834 ;
    wire new_AGEMA_signal_17835 ;
    wire new_AGEMA_signal_17836 ;
    wire new_AGEMA_signal_17837 ;
    wire new_AGEMA_signal_17838 ;
    wire new_AGEMA_signal_17839 ;
    wire new_AGEMA_signal_17840 ;
    wire new_AGEMA_signal_17841 ;
    wire new_AGEMA_signal_17842 ;
    wire new_AGEMA_signal_17843 ;
    wire new_AGEMA_signal_17844 ;
    wire new_AGEMA_signal_17845 ;
    wire new_AGEMA_signal_17846 ;
    wire new_AGEMA_signal_17847 ;
    wire new_AGEMA_signal_17848 ;
    wire new_AGEMA_signal_17849 ;
    wire new_AGEMA_signal_17850 ;
    wire new_AGEMA_signal_17851 ;
    wire new_AGEMA_signal_17852 ;
    wire new_AGEMA_signal_17853 ;
    wire new_AGEMA_signal_17854 ;
    wire new_AGEMA_signal_17855 ;
    wire new_AGEMA_signal_17856 ;
    wire new_AGEMA_signal_17857 ;
    wire new_AGEMA_signal_17858 ;
    wire new_AGEMA_signal_17859 ;
    wire new_AGEMA_signal_17860 ;
    wire new_AGEMA_signal_17861 ;
    wire new_AGEMA_signal_17862 ;
    wire new_AGEMA_signal_17863 ;
    wire new_AGEMA_signal_17864 ;
    wire new_AGEMA_signal_17865 ;
    wire new_AGEMA_signal_17866 ;
    wire new_AGEMA_signal_17867 ;
    wire new_AGEMA_signal_17868 ;
    wire new_AGEMA_signal_17869 ;
    wire new_AGEMA_signal_17870 ;
    wire new_AGEMA_signal_17871 ;
    wire new_AGEMA_signal_17872 ;
    wire new_AGEMA_signal_17873 ;
    wire new_AGEMA_signal_17874 ;
    wire new_AGEMA_signal_17875 ;
    wire new_AGEMA_signal_17876 ;
    wire new_AGEMA_signal_17877 ;
    wire new_AGEMA_signal_17878 ;
    wire new_AGEMA_signal_17879 ;
    wire new_AGEMA_signal_17880 ;
    wire new_AGEMA_signal_17881 ;
    wire new_AGEMA_signal_17882 ;
    wire new_AGEMA_signal_17883 ;
    wire new_AGEMA_signal_17884 ;
    wire new_AGEMA_signal_17885 ;
    wire new_AGEMA_signal_17886 ;
    wire new_AGEMA_signal_17887 ;
    wire new_AGEMA_signal_17888 ;
    wire new_AGEMA_signal_17889 ;
    wire new_AGEMA_signal_17890 ;
    wire new_AGEMA_signal_17891 ;
    wire new_AGEMA_signal_17892 ;
    wire new_AGEMA_signal_17893 ;
    wire new_AGEMA_signal_17894 ;
    wire new_AGEMA_signal_17895 ;
    wire new_AGEMA_signal_17896 ;
    wire new_AGEMA_signal_17897 ;
    wire new_AGEMA_signal_17898 ;
    wire new_AGEMA_signal_17899 ;
    wire new_AGEMA_signal_17900 ;
    wire new_AGEMA_signal_17901 ;
    wire new_AGEMA_signal_17902 ;
    wire new_AGEMA_signal_17903 ;
    wire new_AGEMA_signal_17904 ;
    wire new_AGEMA_signal_17905 ;
    wire new_AGEMA_signal_17906 ;
    wire new_AGEMA_signal_17907 ;
    wire new_AGEMA_signal_17908 ;
    wire new_AGEMA_signal_17909 ;
    wire new_AGEMA_signal_17910 ;
    wire new_AGEMA_signal_17911 ;
    wire new_AGEMA_signal_17912 ;
    wire new_AGEMA_signal_17913 ;
    wire new_AGEMA_signal_17914 ;
    wire new_AGEMA_signal_17915 ;
    wire new_AGEMA_signal_17916 ;
    wire new_AGEMA_signal_17917 ;
    wire new_AGEMA_signal_17918 ;
    wire new_AGEMA_signal_17919 ;
    wire new_AGEMA_signal_17920 ;
    wire new_AGEMA_signal_17921 ;
    wire new_AGEMA_signal_17922 ;
    wire new_AGEMA_signal_17923 ;
    wire new_AGEMA_signal_17924 ;
    wire new_AGEMA_signal_17925 ;
    wire new_AGEMA_signal_17926 ;
    wire new_AGEMA_signal_17927 ;
    wire new_AGEMA_signal_17928 ;
    wire new_AGEMA_signal_17929 ;
    wire new_AGEMA_signal_17930 ;
    wire new_AGEMA_signal_17931 ;
    wire new_AGEMA_signal_17932 ;
    wire new_AGEMA_signal_17933 ;
    wire new_AGEMA_signal_17934 ;
    wire new_AGEMA_signal_17935 ;
    wire new_AGEMA_signal_17936 ;
    wire new_AGEMA_signal_17937 ;
    wire new_AGEMA_signal_17938 ;
    wire new_AGEMA_signal_17939 ;
    wire new_AGEMA_signal_17940 ;
    wire new_AGEMA_signal_17941 ;
    wire new_AGEMA_signal_17942 ;
    wire new_AGEMA_signal_17943 ;
    wire new_AGEMA_signal_17944 ;
    wire new_AGEMA_signal_17945 ;
    wire new_AGEMA_signal_17946 ;
    wire new_AGEMA_signal_17947 ;
    wire new_AGEMA_signal_17948 ;
    wire new_AGEMA_signal_17949 ;
    wire new_AGEMA_signal_17950 ;
    wire new_AGEMA_signal_17951 ;
    wire new_AGEMA_signal_17952 ;
    wire new_AGEMA_signal_17953 ;
    wire new_AGEMA_signal_17954 ;
    wire new_AGEMA_signal_17955 ;
    wire new_AGEMA_signal_17956 ;
    wire new_AGEMA_signal_17957 ;
    wire new_AGEMA_signal_17958 ;
    wire new_AGEMA_signal_17959 ;
    wire new_AGEMA_signal_17960 ;
    wire new_AGEMA_signal_17961 ;
    wire new_AGEMA_signal_17962 ;
    wire new_AGEMA_signal_17963 ;
    wire new_AGEMA_signal_17964 ;
    wire new_AGEMA_signal_17965 ;
    wire new_AGEMA_signal_17966 ;
    wire new_AGEMA_signal_17967 ;
    wire new_AGEMA_signal_17968 ;
    wire new_AGEMA_signal_17969 ;
    wire new_AGEMA_signal_17970 ;
    wire new_AGEMA_signal_17971 ;
    wire new_AGEMA_signal_17972 ;
    wire new_AGEMA_signal_17973 ;
    wire new_AGEMA_signal_17974 ;
    wire new_AGEMA_signal_17975 ;
    wire new_AGEMA_signal_17976 ;
    wire new_AGEMA_signal_17977 ;
    wire new_AGEMA_signal_17978 ;
    wire new_AGEMA_signal_17979 ;
    wire new_AGEMA_signal_17980 ;
    wire new_AGEMA_signal_17981 ;
    wire new_AGEMA_signal_17982 ;
    wire new_AGEMA_signal_17983 ;
    wire new_AGEMA_signal_17984 ;
    wire new_AGEMA_signal_17985 ;
    wire new_AGEMA_signal_17986 ;
    wire new_AGEMA_signal_17987 ;
    wire new_AGEMA_signal_17988 ;
    wire new_AGEMA_signal_17989 ;
    wire new_AGEMA_signal_17990 ;
    wire new_AGEMA_signal_17991 ;
    wire new_AGEMA_signal_17992 ;
    wire new_AGEMA_signal_17993 ;
    wire new_AGEMA_signal_17994 ;
    wire new_AGEMA_signal_17995 ;
    wire new_AGEMA_signal_17996 ;
    wire new_AGEMA_signal_17997 ;
    wire new_AGEMA_signal_17998 ;
    wire new_AGEMA_signal_17999 ;
    wire new_AGEMA_signal_18000 ;
    wire new_AGEMA_signal_18001 ;
    wire new_AGEMA_signal_18002 ;
    wire new_AGEMA_signal_18003 ;
    wire new_AGEMA_signal_18004 ;
    wire new_AGEMA_signal_18005 ;
    wire new_AGEMA_signal_18006 ;
    wire new_AGEMA_signal_18007 ;
    wire new_AGEMA_signal_18008 ;
    wire new_AGEMA_signal_18009 ;
    wire new_AGEMA_signal_18010 ;
    wire new_AGEMA_signal_18011 ;
    wire new_AGEMA_signal_18012 ;
    wire new_AGEMA_signal_18013 ;
    wire new_AGEMA_signal_18014 ;
    wire new_AGEMA_signal_18015 ;
    wire new_AGEMA_signal_18016 ;
    wire new_AGEMA_signal_18017 ;
    wire new_AGEMA_signal_18018 ;
    wire new_AGEMA_signal_18019 ;
    wire new_AGEMA_signal_18020 ;
    wire new_AGEMA_signal_18021 ;
    wire new_AGEMA_signal_18022 ;
    wire new_AGEMA_signal_18023 ;
    wire new_AGEMA_signal_18024 ;
    wire new_AGEMA_signal_18025 ;
    wire new_AGEMA_signal_18026 ;
    wire new_AGEMA_signal_18027 ;
    wire new_AGEMA_signal_18028 ;
    wire new_AGEMA_signal_18029 ;
    wire new_AGEMA_signal_18030 ;
    wire new_AGEMA_signal_18031 ;
    wire new_AGEMA_signal_18032 ;
    wire new_AGEMA_signal_18033 ;
    wire new_AGEMA_signal_18034 ;
    wire new_AGEMA_signal_18035 ;
    wire new_AGEMA_signal_18036 ;
    wire new_AGEMA_signal_18037 ;
    wire new_AGEMA_signal_18038 ;
    wire new_AGEMA_signal_18039 ;
    wire new_AGEMA_signal_18040 ;
    wire new_AGEMA_signal_18041 ;
    wire new_AGEMA_signal_18042 ;
    wire new_AGEMA_signal_18043 ;
    wire new_AGEMA_signal_18044 ;
    wire new_AGEMA_signal_18045 ;
    wire new_AGEMA_signal_18046 ;
    wire new_AGEMA_signal_18047 ;
    wire new_AGEMA_signal_18048 ;
    wire new_AGEMA_signal_18049 ;
    wire new_AGEMA_signal_18050 ;
    wire new_AGEMA_signal_18051 ;
    wire new_AGEMA_signal_18052 ;
    wire new_AGEMA_signal_18053 ;
    wire new_AGEMA_signal_18054 ;
    wire new_AGEMA_signal_18055 ;
    wire new_AGEMA_signal_18056 ;
    wire new_AGEMA_signal_18057 ;
    wire new_AGEMA_signal_18058 ;
    wire new_AGEMA_signal_18059 ;
    wire new_AGEMA_signal_18060 ;
    wire new_AGEMA_signal_18061 ;
    wire new_AGEMA_signal_18062 ;
    wire new_AGEMA_signal_18063 ;
    wire new_AGEMA_signal_18064 ;
    wire new_AGEMA_signal_18065 ;
    wire new_AGEMA_signal_18066 ;
    wire new_AGEMA_signal_18067 ;
    wire new_AGEMA_signal_18068 ;
    wire new_AGEMA_signal_18069 ;
    wire new_AGEMA_signal_18070 ;
    wire new_AGEMA_signal_18071 ;
    wire new_AGEMA_signal_18072 ;
    wire new_AGEMA_signal_18073 ;
    wire new_AGEMA_signal_18074 ;
    wire new_AGEMA_signal_18075 ;
    wire new_AGEMA_signal_18076 ;
    wire new_AGEMA_signal_18077 ;
    wire new_AGEMA_signal_18078 ;
    wire new_AGEMA_signal_18079 ;
    wire new_AGEMA_signal_18080 ;
    wire new_AGEMA_signal_18081 ;
    wire new_AGEMA_signal_18082 ;
    wire new_AGEMA_signal_18083 ;
    wire new_AGEMA_signal_18084 ;
    wire new_AGEMA_signal_18085 ;
    wire new_AGEMA_signal_18086 ;
    wire new_AGEMA_signal_18087 ;
    wire new_AGEMA_signal_18088 ;
    wire new_AGEMA_signal_18089 ;
    wire new_AGEMA_signal_18090 ;
    wire new_AGEMA_signal_18091 ;
    wire new_AGEMA_signal_18092 ;
    wire new_AGEMA_signal_18093 ;
    wire new_AGEMA_signal_18094 ;
    wire new_AGEMA_signal_18095 ;
    wire new_AGEMA_signal_18096 ;
    wire new_AGEMA_signal_18097 ;
    wire new_AGEMA_signal_18098 ;
    wire new_AGEMA_signal_18099 ;
    wire new_AGEMA_signal_18100 ;
    wire new_AGEMA_signal_18101 ;
    wire new_AGEMA_signal_18102 ;
    wire new_AGEMA_signal_18103 ;
    wire new_AGEMA_signal_18104 ;
    wire new_AGEMA_signal_18105 ;
    wire new_AGEMA_signal_18106 ;
    wire new_AGEMA_signal_18107 ;
    wire new_AGEMA_signal_18108 ;
    wire new_AGEMA_signal_18109 ;
    wire new_AGEMA_signal_18110 ;
    wire new_AGEMA_signal_18111 ;
    wire new_AGEMA_signal_18112 ;
    wire new_AGEMA_signal_18113 ;
    wire new_AGEMA_signal_18114 ;
    wire new_AGEMA_signal_18115 ;
    wire new_AGEMA_signal_18116 ;
    wire new_AGEMA_signal_18117 ;
    wire new_AGEMA_signal_18118 ;
    wire new_AGEMA_signal_18119 ;
    wire new_AGEMA_signal_18120 ;
    wire new_AGEMA_signal_18121 ;
    wire new_AGEMA_signal_18122 ;
    wire new_AGEMA_signal_18123 ;
    wire new_AGEMA_signal_18124 ;
    wire new_AGEMA_signal_18125 ;
    wire new_AGEMA_signal_18126 ;
    wire new_AGEMA_signal_18127 ;
    wire new_AGEMA_signal_18128 ;
    wire new_AGEMA_signal_18129 ;
    wire new_AGEMA_signal_18130 ;
    wire new_AGEMA_signal_18131 ;
    wire new_AGEMA_signal_18132 ;
    wire new_AGEMA_signal_18133 ;
    wire new_AGEMA_signal_18134 ;
    wire new_AGEMA_signal_18135 ;
    wire new_AGEMA_signal_18136 ;
    wire new_AGEMA_signal_18137 ;
    wire new_AGEMA_signal_18138 ;
    wire new_AGEMA_signal_18139 ;
    wire new_AGEMA_signal_18140 ;
    wire new_AGEMA_signal_18141 ;
    wire new_AGEMA_signal_18142 ;
    wire new_AGEMA_signal_18143 ;
    wire new_AGEMA_signal_18144 ;
    wire new_AGEMA_signal_18145 ;
    wire new_AGEMA_signal_18146 ;
    wire new_AGEMA_signal_18147 ;
    wire new_AGEMA_signal_18148 ;
    wire new_AGEMA_signal_18149 ;
    wire new_AGEMA_signal_18150 ;
    wire new_AGEMA_signal_18151 ;
    wire new_AGEMA_signal_18152 ;
    wire new_AGEMA_signal_18153 ;
    wire new_AGEMA_signal_18154 ;
    wire new_AGEMA_signal_18155 ;
    wire new_AGEMA_signal_18156 ;
    wire new_AGEMA_signal_18157 ;
    wire new_AGEMA_signal_18158 ;
    wire new_AGEMA_signal_18159 ;
    wire new_AGEMA_signal_18160 ;
    wire new_AGEMA_signal_18161 ;
    wire new_AGEMA_signal_18162 ;
    wire new_AGEMA_signal_18163 ;
    wire new_AGEMA_signal_18164 ;
    wire new_AGEMA_signal_18165 ;
    wire new_AGEMA_signal_18166 ;
    wire new_AGEMA_signal_18167 ;
    wire new_AGEMA_signal_18168 ;
    wire new_AGEMA_signal_18169 ;
    wire new_AGEMA_signal_18170 ;
    wire new_AGEMA_signal_18171 ;
    wire new_AGEMA_signal_18172 ;
    wire new_AGEMA_signal_18173 ;
    wire new_AGEMA_signal_18174 ;
    wire new_AGEMA_signal_18175 ;
    wire new_AGEMA_signal_18176 ;
    wire new_AGEMA_signal_18177 ;
    wire new_AGEMA_signal_18178 ;
    wire new_AGEMA_signal_18179 ;
    wire new_AGEMA_signal_18180 ;
    wire new_AGEMA_signal_18181 ;
    wire new_AGEMA_signal_18182 ;
    wire new_AGEMA_signal_18183 ;
    wire new_AGEMA_signal_18184 ;
    wire new_AGEMA_signal_18185 ;
    wire new_AGEMA_signal_18186 ;
    wire new_AGEMA_signal_18187 ;
    wire new_AGEMA_signal_18188 ;
    wire new_AGEMA_signal_18189 ;
    wire new_AGEMA_signal_18190 ;
    wire new_AGEMA_signal_18191 ;
    wire new_AGEMA_signal_18192 ;
    wire new_AGEMA_signal_18193 ;
    wire new_AGEMA_signal_18194 ;
    wire new_AGEMA_signal_18195 ;
    wire new_AGEMA_signal_18196 ;
    wire new_AGEMA_signal_18197 ;
    wire new_AGEMA_signal_18198 ;
    wire new_AGEMA_signal_18199 ;
    wire new_AGEMA_signal_18200 ;
    wire new_AGEMA_signal_18201 ;
    wire new_AGEMA_signal_18202 ;
    wire new_AGEMA_signal_18203 ;
    wire new_AGEMA_signal_18204 ;
    wire new_AGEMA_signal_18205 ;
    wire new_AGEMA_signal_18206 ;
    wire new_AGEMA_signal_18207 ;
    wire new_AGEMA_signal_18208 ;
    wire new_AGEMA_signal_18209 ;
    wire new_AGEMA_signal_18210 ;
    wire new_AGEMA_signal_18211 ;
    wire new_AGEMA_signal_18212 ;
    wire new_AGEMA_signal_18213 ;
    wire new_AGEMA_signal_18214 ;
    wire new_AGEMA_signal_18215 ;
    wire new_AGEMA_signal_18216 ;
    wire new_AGEMA_signal_18217 ;
    wire new_AGEMA_signal_18218 ;
    wire new_AGEMA_signal_18219 ;
    wire new_AGEMA_signal_18220 ;
    wire new_AGEMA_signal_18221 ;
    wire new_AGEMA_signal_18222 ;
    wire new_AGEMA_signal_18223 ;
    wire new_AGEMA_signal_18224 ;
    wire new_AGEMA_signal_18225 ;
    wire new_AGEMA_signal_18226 ;
    wire new_AGEMA_signal_18227 ;
    wire new_AGEMA_signal_18228 ;
    wire new_AGEMA_signal_18229 ;
    wire new_AGEMA_signal_18230 ;
    wire new_AGEMA_signal_18231 ;
    wire new_AGEMA_signal_18232 ;
    wire new_AGEMA_signal_18233 ;
    wire new_AGEMA_signal_18234 ;
    wire new_AGEMA_signal_18235 ;
    wire new_AGEMA_signal_18236 ;
    wire new_AGEMA_signal_18237 ;
    wire new_AGEMA_signal_18238 ;
    wire new_AGEMA_signal_18239 ;
    wire new_AGEMA_signal_18240 ;
    wire new_AGEMA_signal_18241 ;
    wire new_AGEMA_signal_18242 ;
    wire new_AGEMA_signal_18243 ;
    wire new_AGEMA_signal_18244 ;
    wire new_AGEMA_signal_18245 ;
    wire new_AGEMA_signal_18246 ;
    wire new_AGEMA_signal_18247 ;
    wire new_AGEMA_signal_18248 ;
    wire new_AGEMA_signal_18249 ;
    wire new_AGEMA_signal_18250 ;
    wire new_AGEMA_signal_18251 ;
    wire new_AGEMA_signal_18252 ;
    wire new_AGEMA_signal_18253 ;
    wire new_AGEMA_signal_18254 ;
    wire new_AGEMA_signal_18255 ;
    wire new_AGEMA_signal_18256 ;
    wire new_AGEMA_signal_18257 ;
    wire new_AGEMA_signal_18258 ;
    wire new_AGEMA_signal_18259 ;
    wire new_AGEMA_signal_18260 ;
    wire new_AGEMA_signal_18261 ;
    wire new_AGEMA_signal_18262 ;
    wire new_AGEMA_signal_18263 ;
    wire new_AGEMA_signal_18264 ;
    wire new_AGEMA_signal_18265 ;
    wire new_AGEMA_signal_18266 ;
    wire new_AGEMA_signal_18267 ;
    wire new_AGEMA_signal_18268 ;
    wire new_AGEMA_signal_18269 ;
    wire new_AGEMA_signal_18270 ;
    wire new_AGEMA_signal_18271 ;
    wire new_AGEMA_signal_18272 ;
    wire new_AGEMA_signal_18273 ;
    wire new_AGEMA_signal_18274 ;
    wire new_AGEMA_signal_18275 ;
    wire new_AGEMA_signal_18276 ;
    wire new_AGEMA_signal_18277 ;
    wire new_AGEMA_signal_18278 ;
    wire new_AGEMA_signal_18279 ;
    wire new_AGEMA_signal_18280 ;
    wire new_AGEMA_signal_18281 ;
    wire new_AGEMA_signal_18282 ;
    wire new_AGEMA_signal_18283 ;
    wire new_AGEMA_signal_18284 ;
    wire new_AGEMA_signal_18285 ;
    wire new_AGEMA_signal_18286 ;
    wire new_AGEMA_signal_18287 ;
    wire new_AGEMA_signal_18288 ;
    wire new_AGEMA_signal_18289 ;
    wire new_AGEMA_signal_18290 ;
    wire new_AGEMA_signal_18291 ;
    wire new_AGEMA_signal_18292 ;
    wire new_AGEMA_signal_18293 ;
    wire new_AGEMA_signal_18294 ;
    wire new_AGEMA_signal_18295 ;
    wire new_AGEMA_signal_18296 ;
    wire new_AGEMA_signal_18297 ;
    wire new_AGEMA_signal_18298 ;
    wire new_AGEMA_signal_18299 ;
    wire new_AGEMA_signal_18300 ;
    wire new_AGEMA_signal_18301 ;
    wire new_AGEMA_signal_18302 ;
    wire new_AGEMA_signal_18303 ;
    wire new_AGEMA_signal_18304 ;
    wire new_AGEMA_signal_18305 ;
    wire new_AGEMA_signal_18306 ;
    wire new_AGEMA_signal_18307 ;
    wire new_AGEMA_signal_18308 ;
    wire new_AGEMA_signal_18309 ;
    wire new_AGEMA_signal_18310 ;
    wire new_AGEMA_signal_18311 ;
    wire new_AGEMA_signal_18312 ;
    wire new_AGEMA_signal_18313 ;
    wire new_AGEMA_signal_18314 ;
    wire new_AGEMA_signal_18315 ;
    wire new_AGEMA_signal_18316 ;
    wire new_AGEMA_signal_18317 ;
    wire new_AGEMA_signal_18318 ;
    wire new_AGEMA_signal_18319 ;
    wire new_AGEMA_signal_18320 ;
    wire new_AGEMA_signal_18321 ;
    wire new_AGEMA_signal_18322 ;
    wire new_AGEMA_signal_18323 ;
    wire new_AGEMA_signal_18324 ;
    wire new_AGEMA_signal_18325 ;
    wire new_AGEMA_signal_18326 ;
    wire new_AGEMA_signal_18327 ;
    wire new_AGEMA_signal_18328 ;
    wire new_AGEMA_signal_18329 ;
    wire new_AGEMA_signal_18330 ;
    wire new_AGEMA_signal_18331 ;
    wire new_AGEMA_signal_18332 ;
    wire new_AGEMA_signal_18333 ;
    wire new_AGEMA_signal_18334 ;
    wire new_AGEMA_signal_18335 ;
    wire new_AGEMA_signal_18336 ;
    wire new_AGEMA_signal_18337 ;
    wire new_AGEMA_signal_18338 ;
    wire new_AGEMA_signal_18339 ;
    wire new_AGEMA_signal_18340 ;
    wire new_AGEMA_signal_18341 ;
    wire new_AGEMA_signal_18342 ;
    wire new_AGEMA_signal_18343 ;
    wire new_AGEMA_signal_18344 ;
    wire new_AGEMA_signal_18345 ;
    wire new_AGEMA_signal_18346 ;
    wire new_AGEMA_signal_18347 ;
    wire new_AGEMA_signal_18348 ;
    wire new_AGEMA_signal_18349 ;
    wire new_AGEMA_signal_18350 ;
    wire new_AGEMA_signal_18351 ;
    wire new_AGEMA_signal_18352 ;
    wire new_AGEMA_signal_18353 ;
    wire new_AGEMA_signal_18354 ;
    wire new_AGEMA_signal_18355 ;
    wire new_AGEMA_signal_18356 ;
    wire new_AGEMA_signal_18357 ;
    wire new_AGEMA_signal_18358 ;
    wire new_AGEMA_signal_18359 ;
    wire new_AGEMA_signal_18360 ;
    wire new_AGEMA_signal_18361 ;
    wire new_AGEMA_signal_18362 ;
    wire new_AGEMA_signal_18363 ;
    wire new_AGEMA_signal_18364 ;
    wire new_AGEMA_signal_18365 ;
    wire new_AGEMA_signal_18366 ;
    wire new_AGEMA_signal_18367 ;
    wire new_AGEMA_signal_18368 ;
    wire new_AGEMA_signal_18369 ;
    wire new_AGEMA_signal_18370 ;
    wire new_AGEMA_signal_18371 ;
    wire new_AGEMA_signal_18372 ;
    wire new_AGEMA_signal_18373 ;
    wire new_AGEMA_signal_18374 ;
    wire new_AGEMA_signal_18375 ;
    wire new_AGEMA_signal_18376 ;
    wire new_AGEMA_signal_18377 ;
    wire new_AGEMA_signal_18378 ;
    wire new_AGEMA_signal_18379 ;
    wire new_AGEMA_signal_18380 ;
    wire new_AGEMA_signal_18381 ;
    wire new_AGEMA_signal_18382 ;
    wire new_AGEMA_signal_18383 ;
    wire new_AGEMA_signal_18384 ;
    wire new_AGEMA_signal_18385 ;
    wire new_AGEMA_signal_18386 ;
    wire new_AGEMA_signal_18387 ;
    wire new_AGEMA_signal_18388 ;
    wire new_AGEMA_signal_18389 ;
    wire new_AGEMA_signal_18390 ;
    wire new_AGEMA_signal_18391 ;
    wire new_AGEMA_signal_18392 ;
    wire new_AGEMA_signal_18393 ;
    wire new_AGEMA_signal_18394 ;
    wire new_AGEMA_signal_18395 ;
    wire new_AGEMA_signal_18396 ;
    wire new_AGEMA_signal_18397 ;
    wire new_AGEMA_signal_18398 ;
    wire new_AGEMA_signal_18399 ;
    wire new_AGEMA_signal_18400 ;
    wire new_AGEMA_signal_18401 ;
    wire new_AGEMA_signal_18402 ;
    wire new_AGEMA_signal_18403 ;
    wire new_AGEMA_signal_18404 ;
    wire new_AGEMA_signal_18405 ;
    wire new_AGEMA_signal_18406 ;
    wire new_AGEMA_signal_18407 ;
    wire new_AGEMA_signal_18408 ;
    wire new_AGEMA_signal_18409 ;
    wire new_AGEMA_signal_18410 ;
    wire new_AGEMA_signal_18411 ;
    wire new_AGEMA_signal_18412 ;
    wire new_AGEMA_signal_18413 ;
    wire new_AGEMA_signal_18414 ;
    wire new_AGEMA_signal_18415 ;
    wire new_AGEMA_signal_18416 ;
    wire new_AGEMA_signal_18417 ;
    wire new_AGEMA_signal_18418 ;
    wire new_AGEMA_signal_18419 ;
    wire new_AGEMA_signal_18420 ;
    wire new_AGEMA_signal_18421 ;
    wire new_AGEMA_signal_18422 ;
    wire new_AGEMA_signal_18423 ;
    wire new_AGEMA_signal_18424 ;
    wire new_AGEMA_signal_18425 ;
    wire new_AGEMA_signal_18426 ;
    wire new_AGEMA_signal_18427 ;
    wire new_AGEMA_signal_18428 ;
    wire new_AGEMA_signal_18429 ;
    wire new_AGEMA_signal_18430 ;
    wire new_AGEMA_signal_18431 ;
    wire new_AGEMA_signal_18432 ;
    wire new_AGEMA_signal_18433 ;
    wire new_AGEMA_signal_18434 ;
    wire new_AGEMA_signal_18435 ;
    wire new_AGEMA_signal_18436 ;
    wire new_AGEMA_signal_18437 ;
    wire new_AGEMA_signal_18438 ;
    wire new_AGEMA_signal_18439 ;
    wire new_AGEMA_signal_18440 ;
    wire new_AGEMA_signal_18441 ;
    wire new_AGEMA_signal_18442 ;
    wire new_AGEMA_signal_18443 ;
    wire new_AGEMA_signal_18444 ;
    wire new_AGEMA_signal_18445 ;
    wire new_AGEMA_signal_18446 ;
    wire new_AGEMA_signal_18447 ;
    wire new_AGEMA_signal_18448 ;
    wire new_AGEMA_signal_18449 ;
    wire new_AGEMA_signal_18450 ;
    wire new_AGEMA_signal_18451 ;
    wire new_AGEMA_signal_18452 ;
    wire new_AGEMA_signal_18453 ;
    wire new_AGEMA_signal_18454 ;
    wire new_AGEMA_signal_18455 ;
    wire new_AGEMA_signal_18456 ;
    wire new_AGEMA_signal_18457 ;
    wire new_AGEMA_signal_18458 ;
    wire new_AGEMA_signal_18459 ;
    wire new_AGEMA_signal_18460 ;
    wire new_AGEMA_signal_18461 ;
    wire new_AGEMA_signal_18462 ;
    wire new_AGEMA_signal_18463 ;
    wire new_AGEMA_signal_18464 ;
    wire new_AGEMA_signal_18465 ;
    wire new_AGEMA_signal_18466 ;
    wire new_AGEMA_signal_18467 ;
    wire new_AGEMA_signal_18468 ;
    wire new_AGEMA_signal_18469 ;
    wire new_AGEMA_signal_18470 ;
    wire new_AGEMA_signal_18471 ;
    wire new_AGEMA_signal_18472 ;
    wire new_AGEMA_signal_18473 ;
    wire new_AGEMA_signal_18474 ;
    wire new_AGEMA_signal_18475 ;
    wire new_AGEMA_signal_18476 ;
    wire new_AGEMA_signal_18477 ;
    wire new_AGEMA_signal_18478 ;
    wire new_AGEMA_signal_18479 ;
    wire new_AGEMA_signal_18480 ;
    wire new_AGEMA_signal_18481 ;
    wire new_AGEMA_signal_18482 ;
    wire new_AGEMA_signal_18483 ;
    wire new_AGEMA_signal_18484 ;
    wire new_AGEMA_signal_18485 ;
    wire new_AGEMA_signal_18486 ;
    wire new_AGEMA_signal_18487 ;
    wire new_AGEMA_signal_18488 ;
    wire new_AGEMA_signal_18489 ;
    wire new_AGEMA_signal_18490 ;
    wire new_AGEMA_signal_18491 ;
    wire new_AGEMA_signal_18492 ;
    wire new_AGEMA_signal_18493 ;
    wire new_AGEMA_signal_18494 ;
    wire new_AGEMA_signal_18495 ;
    wire new_AGEMA_signal_18496 ;
    wire new_AGEMA_signal_18497 ;
    wire new_AGEMA_signal_18498 ;
    wire new_AGEMA_signal_18499 ;
    wire new_AGEMA_signal_18500 ;
    wire new_AGEMA_signal_18501 ;
    wire new_AGEMA_signal_18502 ;
    wire new_AGEMA_signal_18503 ;
    wire new_AGEMA_signal_18504 ;
    wire new_AGEMA_signal_18505 ;
    wire new_AGEMA_signal_18506 ;
    wire new_AGEMA_signal_18507 ;
    wire new_AGEMA_signal_18508 ;
    wire new_AGEMA_signal_18509 ;
    wire new_AGEMA_signal_18510 ;
    wire new_AGEMA_signal_18511 ;
    wire new_AGEMA_signal_18512 ;
    wire new_AGEMA_signal_18513 ;
    wire new_AGEMA_signal_18514 ;
    wire new_AGEMA_signal_18515 ;
    wire new_AGEMA_signal_18516 ;
    wire new_AGEMA_signal_18517 ;
    wire new_AGEMA_signal_18518 ;
    wire new_AGEMA_signal_18519 ;
    wire new_AGEMA_signal_18520 ;
    wire new_AGEMA_signal_18521 ;
    wire new_AGEMA_signal_18522 ;
    wire new_AGEMA_signal_18523 ;
    wire new_AGEMA_signal_18524 ;
    wire new_AGEMA_signal_18525 ;
    wire new_AGEMA_signal_18526 ;
    wire new_AGEMA_signal_18527 ;
    wire new_AGEMA_signal_18528 ;
    wire new_AGEMA_signal_18529 ;
    wire new_AGEMA_signal_18530 ;
    wire new_AGEMA_signal_18531 ;
    wire new_AGEMA_signal_18532 ;
    wire new_AGEMA_signal_18533 ;
    wire new_AGEMA_signal_18534 ;
    wire new_AGEMA_signal_18535 ;
    wire new_AGEMA_signal_18536 ;
    wire new_AGEMA_signal_18537 ;
    wire new_AGEMA_signal_18538 ;
    wire new_AGEMA_signal_18539 ;
    wire new_AGEMA_signal_18540 ;
    wire new_AGEMA_signal_18541 ;
    wire new_AGEMA_signal_18542 ;
    wire new_AGEMA_signal_18543 ;
    wire new_AGEMA_signal_18544 ;
    wire new_AGEMA_signal_18545 ;
    wire new_AGEMA_signal_18546 ;
    wire new_AGEMA_signal_18547 ;
    wire new_AGEMA_signal_18548 ;
    wire new_AGEMA_signal_18549 ;
    wire new_AGEMA_signal_18550 ;
    wire new_AGEMA_signal_18551 ;
    wire new_AGEMA_signal_18552 ;
    wire new_AGEMA_signal_18553 ;
    wire new_AGEMA_signal_18554 ;
    wire new_AGEMA_signal_18555 ;
    wire new_AGEMA_signal_18556 ;
    wire new_AGEMA_signal_18557 ;
    wire new_AGEMA_signal_18558 ;
    wire new_AGEMA_signal_18559 ;
    wire new_AGEMA_signal_18560 ;
    wire new_AGEMA_signal_18561 ;
    wire new_AGEMA_signal_18562 ;
    wire new_AGEMA_signal_18563 ;
    wire new_AGEMA_signal_18564 ;
    wire new_AGEMA_signal_18565 ;
    wire new_AGEMA_signal_18566 ;
    wire new_AGEMA_signal_18567 ;
    wire new_AGEMA_signal_18568 ;
    wire new_AGEMA_signal_18569 ;
    wire new_AGEMA_signal_18570 ;
    wire new_AGEMA_signal_18571 ;
    wire new_AGEMA_signal_18572 ;
    wire new_AGEMA_signal_18573 ;
    wire new_AGEMA_signal_18574 ;
    wire new_AGEMA_signal_18575 ;
    wire new_AGEMA_signal_18576 ;
    wire new_AGEMA_signal_18577 ;
    wire new_AGEMA_signal_18578 ;
    wire new_AGEMA_signal_18579 ;
    wire new_AGEMA_signal_18580 ;
    wire new_AGEMA_signal_18581 ;
    wire new_AGEMA_signal_18582 ;
    wire new_AGEMA_signal_18583 ;
    wire new_AGEMA_signal_18584 ;
    wire new_AGEMA_signal_18585 ;
    wire new_AGEMA_signal_18586 ;
    wire new_AGEMA_signal_18587 ;
    wire new_AGEMA_signal_18588 ;
    wire new_AGEMA_signal_18589 ;
    wire new_AGEMA_signal_18590 ;
    wire new_AGEMA_signal_18591 ;
    wire new_AGEMA_signal_18592 ;
    wire new_AGEMA_signal_18593 ;
    wire new_AGEMA_signal_18594 ;
    wire new_AGEMA_signal_18595 ;
    wire new_AGEMA_signal_18596 ;
    wire new_AGEMA_signal_18597 ;
    wire new_AGEMA_signal_18598 ;
    wire new_AGEMA_signal_18599 ;
    wire new_AGEMA_signal_18600 ;
    wire new_AGEMA_signal_18601 ;
    wire new_AGEMA_signal_18602 ;
    wire new_AGEMA_signal_18603 ;
    wire new_AGEMA_signal_18604 ;
    wire new_AGEMA_signal_18605 ;
    wire new_AGEMA_signal_18606 ;
    wire new_AGEMA_signal_18607 ;
    wire new_AGEMA_signal_18608 ;
    wire new_AGEMA_signal_18609 ;
    wire new_AGEMA_signal_18610 ;
    wire new_AGEMA_signal_18611 ;
    wire new_AGEMA_signal_18612 ;
    wire new_AGEMA_signal_18613 ;
    wire new_AGEMA_signal_18614 ;
    wire new_AGEMA_signal_18615 ;
    wire new_AGEMA_signal_18616 ;
    wire new_AGEMA_signal_18617 ;
    wire new_AGEMA_signal_18618 ;
    wire new_AGEMA_signal_18619 ;
    wire new_AGEMA_signal_18620 ;
    wire new_AGEMA_signal_18621 ;
    wire new_AGEMA_signal_18622 ;
    wire new_AGEMA_signal_18623 ;
    wire new_AGEMA_signal_18624 ;
    wire new_AGEMA_signal_18625 ;
    wire new_AGEMA_signal_18626 ;
    wire new_AGEMA_signal_18627 ;
    wire new_AGEMA_signal_18628 ;
    wire new_AGEMA_signal_18629 ;
    wire new_AGEMA_signal_18630 ;
    wire new_AGEMA_signal_18631 ;
    wire new_AGEMA_signal_18632 ;
    wire new_AGEMA_signal_18633 ;
    wire new_AGEMA_signal_18634 ;
    wire new_AGEMA_signal_18635 ;
    wire new_AGEMA_signal_18636 ;
    wire new_AGEMA_signal_18637 ;
    wire new_AGEMA_signal_18638 ;
    wire new_AGEMA_signal_18639 ;
    wire new_AGEMA_signal_18640 ;
    wire new_AGEMA_signal_18641 ;
    wire new_AGEMA_signal_18642 ;
    wire new_AGEMA_signal_18643 ;
    wire new_AGEMA_signal_18644 ;
    wire new_AGEMA_signal_18645 ;
    wire new_AGEMA_signal_18646 ;
    wire new_AGEMA_signal_18647 ;
    wire new_AGEMA_signal_18648 ;
    wire new_AGEMA_signal_18649 ;
    wire new_AGEMA_signal_18650 ;
    wire new_AGEMA_signal_18651 ;
    wire new_AGEMA_signal_18652 ;
    wire new_AGEMA_signal_18653 ;
    wire new_AGEMA_signal_18654 ;
    wire new_AGEMA_signal_18655 ;
    wire new_AGEMA_signal_18656 ;
    wire new_AGEMA_signal_18657 ;
    wire new_AGEMA_signal_18658 ;
    wire new_AGEMA_signal_18659 ;
    wire new_AGEMA_signal_18660 ;
    wire new_AGEMA_signal_18661 ;
    wire new_AGEMA_signal_18662 ;
    wire new_AGEMA_signal_18663 ;
    wire new_AGEMA_signal_18664 ;
    wire new_AGEMA_signal_18665 ;
    wire new_AGEMA_signal_18666 ;
    wire new_AGEMA_signal_18667 ;
    wire new_AGEMA_signal_18668 ;
    wire new_AGEMA_signal_18669 ;
    wire new_AGEMA_signal_18670 ;
    wire new_AGEMA_signal_18671 ;
    wire new_AGEMA_signal_18672 ;
    wire new_AGEMA_signal_18673 ;
    wire new_AGEMA_signal_18674 ;
    wire new_AGEMA_signal_18675 ;
    wire new_AGEMA_signal_18676 ;
    wire new_AGEMA_signal_18677 ;
    wire new_AGEMA_signal_18678 ;
    wire new_AGEMA_signal_18679 ;
    wire new_AGEMA_signal_18680 ;
    wire new_AGEMA_signal_18681 ;
    wire new_AGEMA_signal_18682 ;
    wire new_AGEMA_signal_18683 ;
    wire new_AGEMA_signal_18684 ;
    wire new_AGEMA_signal_18685 ;
    wire new_AGEMA_signal_18686 ;
    wire new_AGEMA_signal_18687 ;
    wire new_AGEMA_signal_18688 ;
    wire new_AGEMA_signal_18689 ;
    wire new_AGEMA_signal_18690 ;
    wire new_AGEMA_signal_18691 ;
    wire new_AGEMA_signal_18692 ;
    wire new_AGEMA_signal_18693 ;
    wire new_AGEMA_signal_18694 ;
    wire new_AGEMA_signal_18695 ;
    wire new_AGEMA_signal_18696 ;
    wire new_AGEMA_signal_18697 ;
    wire new_AGEMA_signal_18698 ;
    wire new_AGEMA_signal_18699 ;
    wire new_AGEMA_signal_18700 ;
    wire new_AGEMA_signal_18701 ;
    wire new_AGEMA_signal_18702 ;
    wire new_AGEMA_signal_18703 ;
    wire new_AGEMA_signal_18704 ;
    wire new_AGEMA_signal_18705 ;
    wire new_AGEMA_signal_18706 ;
    wire new_AGEMA_signal_18707 ;
    wire new_AGEMA_signal_18708 ;
    wire new_AGEMA_signal_18709 ;
    wire new_AGEMA_signal_18710 ;
    wire new_AGEMA_signal_18711 ;
    wire new_AGEMA_signal_18712 ;
    wire new_AGEMA_signal_18713 ;
    wire new_AGEMA_signal_18714 ;
    wire new_AGEMA_signal_18715 ;
    wire new_AGEMA_signal_18716 ;
    wire new_AGEMA_signal_18717 ;
    wire new_AGEMA_signal_18718 ;
    wire new_AGEMA_signal_18719 ;
    wire new_AGEMA_signal_18720 ;
    wire new_AGEMA_signal_18721 ;
    wire new_AGEMA_signal_18722 ;
    wire new_AGEMA_signal_18723 ;
    wire new_AGEMA_signal_18724 ;
    wire new_AGEMA_signal_18725 ;
    wire new_AGEMA_signal_18726 ;
    wire new_AGEMA_signal_18727 ;
    wire new_AGEMA_signal_18728 ;
    wire new_AGEMA_signal_18729 ;
    wire new_AGEMA_signal_18730 ;
    wire new_AGEMA_signal_18731 ;
    wire new_AGEMA_signal_18732 ;
    wire new_AGEMA_signal_18733 ;
    wire new_AGEMA_signal_18734 ;
    wire new_AGEMA_signal_18735 ;
    wire new_AGEMA_signal_18736 ;
    wire new_AGEMA_signal_18737 ;
    wire new_AGEMA_signal_18738 ;
    wire new_AGEMA_signal_18739 ;
    wire new_AGEMA_signal_18740 ;
    wire new_AGEMA_signal_18741 ;
    wire new_AGEMA_signal_18742 ;
    wire new_AGEMA_signal_18743 ;
    wire new_AGEMA_signal_18744 ;
    wire new_AGEMA_signal_18745 ;
    wire new_AGEMA_signal_18746 ;
    wire new_AGEMA_signal_18747 ;
    wire new_AGEMA_signal_18748 ;
    wire new_AGEMA_signal_18749 ;
    wire new_AGEMA_signal_18750 ;
    wire new_AGEMA_signal_18751 ;
    wire new_AGEMA_signal_18752 ;
    wire new_AGEMA_signal_18753 ;
    wire new_AGEMA_signal_18754 ;
    wire new_AGEMA_signal_18755 ;
    wire new_AGEMA_signal_18756 ;
    wire new_AGEMA_signal_18757 ;
    wire new_AGEMA_signal_18758 ;
    wire new_AGEMA_signal_18759 ;
    wire new_AGEMA_signal_18760 ;
    wire new_AGEMA_signal_18761 ;
    wire new_AGEMA_signal_18762 ;
    wire new_AGEMA_signal_18763 ;
    wire new_AGEMA_signal_18764 ;
    wire new_AGEMA_signal_18765 ;
    wire new_AGEMA_signal_18766 ;
    wire new_AGEMA_signal_18767 ;
    wire new_AGEMA_signal_18768 ;
    wire new_AGEMA_signal_18769 ;
    wire new_AGEMA_signal_18770 ;
    wire new_AGEMA_signal_18771 ;
    wire new_AGEMA_signal_18772 ;
    wire new_AGEMA_signal_18773 ;
    wire new_AGEMA_signal_18774 ;
    wire new_AGEMA_signal_18775 ;
    wire new_AGEMA_signal_18776 ;
    wire new_AGEMA_signal_18777 ;
    wire new_AGEMA_signal_18778 ;
    wire new_AGEMA_signal_18779 ;
    wire new_AGEMA_signal_18780 ;
    wire new_AGEMA_signal_18781 ;
    wire new_AGEMA_signal_18782 ;
    wire new_AGEMA_signal_18783 ;
    wire new_AGEMA_signal_18784 ;
    wire new_AGEMA_signal_18785 ;
    wire new_AGEMA_signal_18786 ;
    wire new_AGEMA_signal_18787 ;
    wire new_AGEMA_signal_18788 ;
    wire new_AGEMA_signal_18789 ;
    wire new_AGEMA_signal_18790 ;
    wire new_AGEMA_signal_18791 ;
    wire new_AGEMA_signal_18792 ;
    wire new_AGEMA_signal_18793 ;
    wire new_AGEMA_signal_18794 ;
    wire new_AGEMA_signal_18795 ;
    wire new_AGEMA_signal_18796 ;
    wire new_AGEMA_signal_18797 ;
    wire new_AGEMA_signal_18798 ;
    wire new_AGEMA_signal_18799 ;
    wire new_AGEMA_signal_18800 ;
    wire new_AGEMA_signal_18801 ;
    wire new_AGEMA_signal_18802 ;
    wire new_AGEMA_signal_18803 ;
    wire new_AGEMA_signal_18804 ;
    wire new_AGEMA_signal_18805 ;
    wire new_AGEMA_signal_18806 ;
    wire new_AGEMA_signal_18807 ;
    wire new_AGEMA_signal_18808 ;
    wire new_AGEMA_signal_18809 ;
    wire new_AGEMA_signal_18810 ;
    wire new_AGEMA_signal_18811 ;
    wire new_AGEMA_signal_18812 ;
    wire new_AGEMA_signal_18813 ;
    wire new_AGEMA_signal_18814 ;
    wire new_AGEMA_signal_18815 ;
    wire new_AGEMA_signal_18816 ;
    wire new_AGEMA_signal_18817 ;
    wire new_AGEMA_signal_18818 ;
    wire new_AGEMA_signal_18819 ;
    wire new_AGEMA_signal_18820 ;
    wire new_AGEMA_signal_18821 ;
    wire new_AGEMA_signal_18822 ;
    wire new_AGEMA_signal_18823 ;
    wire new_AGEMA_signal_18824 ;
    wire new_AGEMA_signal_18825 ;
    wire new_AGEMA_signal_18826 ;
    wire new_AGEMA_signal_18827 ;
    wire new_AGEMA_signal_18828 ;
    wire new_AGEMA_signal_18829 ;
    wire new_AGEMA_signal_18830 ;
    wire new_AGEMA_signal_18831 ;
    wire new_AGEMA_signal_18832 ;
    wire new_AGEMA_signal_18833 ;
    wire new_AGEMA_signal_18834 ;
    wire new_AGEMA_signal_18835 ;
    wire new_AGEMA_signal_18836 ;
    wire new_AGEMA_signal_18837 ;
    wire new_AGEMA_signal_18838 ;
    wire new_AGEMA_signal_18839 ;
    wire new_AGEMA_signal_18840 ;
    wire new_AGEMA_signal_18841 ;
    wire new_AGEMA_signal_18842 ;
    wire new_AGEMA_signal_18843 ;
    wire new_AGEMA_signal_18844 ;
    wire new_AGEMA_signal_18845 ;
    wire new_AGEMA_signal_18846 ;
    wire new_AGEMA_signal_18847 ;
    wire new_AGEMA_signal_18848 ;
    wire new_AGEMA_signal_18849 ;
    wire new_AGEMA_signal_18850 ;
    wire new_AGEMA_signal_18851 ;
    wire new_AGEMA_signal_18852 ;
    wire new_AGEMA_signal_18853 ;
    wire new_AGEMA_signal_18854 ;
    wire new_AGEMA_signal_18855 ;
    wire new_AGEMA_signal_18856 ;
    wire new_AGEMA_signal_18857 ;
    wire new_AGEMA_signal_18858 ;
    wire new_AGEMA_signal_18859 ;
    wire new_AGEMA_signal_18860 ;
    wire new_AGEMA_signal_18861 ;
    wire new_AGEMA_signal_18862 ;
    wire new_AGEMA_signal_18863 ;
    wire new_AGEMA_signal_18864 ;
    wire new_AGEMA_signal_18865 ;
    wire new_AGEMA_signal_18866 ;
    wire new_AGEMA_signal_18867 ;
    wire new_AGEMA_signal_18868 ;
    wire new_AGEMA_signal_18869 ;
    wire new_AGEMA_signal_18870 ;
    wire new_AGEMA_signal_18871 ;
    wire new_AGEMA_signal_18872 ;
    wire new_AGEMA_signal_18873 ;
    wire new_AGEMA_signal_18874 ;
    wire new_AGEMA_signal_18875 ;
    wire new_AGEMA_signal_18876 ;
    wire new_AGEMA_signal_18877 ;
    wire new_AGEMA_signal_18878 ;
    wire new_AGEMA_signal_18879 ;
    wire new_AGEMA_signal_18880 ;
    wire new_AGEMA_signal_18881 ;
    wire new_AGEMA_signal_18882 ;
    wire new_AGEMA_signal_18883 ;
    wire new_AGEMA_signal_18884 ;
    wire new_AGEMA_signal_18885 ;
    wire new_AGEMA_signal_18886 ;
    wire new_AGEMA_signal_18887 ;
    wire new_AGEMA_signal_18888 ;
    wire new_AGEMA_signal_18889 ;
    wire new_AGEMA_signal_18890 ;
    wire new_AGEMA_signal_18891 ;
    wire new_AGEMA_signal_18892 ;
    wire new_AGEMA_signal_18893 ;
    wire new_AGEMA_signal_18894 ;
    wire new_AGEMA_signal_18895 ;
    wire new_AGEMA_signal_18896 ;
    wire new_AGEMA_signal_18897 ;
    wire new_AGEMA_signal_18898 ;
    wire new_AGEMA_signal_18899 ;
    wire new_AGEMA_signal_18900 ;
    wire new_AGEMA_signal_18901 ;
    wire new_AGEMA_signal_18902 ;
    wire new_AGEMA_signal_18903 ;
    wire new_AGEMA_signal_18904 ;
    wire new_AGEMA_signal_18905 ;
    wire new_AGEMA_signal_18906 ;
    wire new_AGEMA_signal_18907 ;
    wire new_AGEMA_signal_18908 ;
    wire new_AGEMA_signal_18909 ;
    wire new_AGEMA_signal_18910 ;
    wire new_AGEMA_signal_18911 ;
    wire new_AGEMA_signal_18912 ;
    wire new_AGEMA_signal_18913 ;
    wire new_AGEMA_signal_18914 ;
    wire new_AGEMA_signal_18915 ;
    wire new_AGEMA_signal_18916 ;
    wire new_AGEMA_signal_18917 ;
    wire new_AGEMA_signal_18918 ;
    wire new_AGEMA_signal_18919 ;
    wire new_AGEMA_signal_18920 ;
    wire new_AGEMA_signal_18921 ;
    wire new_AGEMA_signal_18922 ;
    wire new_AGEMA_signal_18923 ;
    wire new_AGEMA_signal_18924 ;
    wire new_AGEMA_signal_18925 ;
    wire new_AGEMA_signal_18926 ;
    wire new_AGEMA_signal_18927 ;
    wire new_AGEMA_signal_18928 ;
    wire new_AGEMA_signal_18929 ;
    wire new_AGEMA_signal_18930 ;
    wire new_AGEMA_signal_18931 ;
    wire new_AGEMA_signal_18932 ;
    wire new_AGEMA_signal_18933 ;
    wire new_AGEMA_signal_18934 ;
    wire new_AGEMA_signal_18935 ;
    wire new_AGEMA_signal_18936 ;
    wire new_AGEMA_signal_18937 ;
    wire new_AGEMA_signal_18938 ;
    wire new_AGEMA_signal_18939 ;
    wire new_AGEMA_signal_18940 ;
    wire new_AGEMA_signal_18941 ;
    wire new_AGEMA_signal_18942 ;
    wire new_AGEMA_signal_18943 ;
    wire new_AGEMA_signal_18944 ;
    wire new_AGEMA_signal_18945 ;
    wire new_AGEMA_signal_18946 ;
    wire new_AGEMA_signal_18947 ;
    wire new_AGEMA_signal_18948 ;
    wire new_AGEMA_signal_18949 ;
    wire new_AGEMA_signal_18950 ;
    wire new_AGEMA_signal_18951 ;
    wire new_AGEMA_signal_18952 ;
    wire new_AGEMA_signal_18953 ;
    wire new_AGEMA_signal_18954 ;
    wire new_AGEMA_signal_18955 ;
    wire new_AGEMA_signal_18956 ;
    wire new_AGEMA_signal_18957 ;
    wire new_AGEMA_signal_18958 ;
    wire new_AGEMA_signal_18959 ;
    wire new_AGEMA_signal_18960 ;
    wire new_AGEMA_signal_18961 ;
    wire new_AGEMA_signal_18962 ;
    wire new_AGEMA_signal_18963 ;
    wire new_AGEMA_signal_18964 ;
    wire new_AGEMA_signal_18965 ;
    wire new_AGEMA_signal_18966 ;
    wire new_AGEMA_signal_18967 ;
    wire new_AGEMA_signal_18968 ;
    wire new_AGEMA_signal_18969 ;
    wire new_AGEMA_signal_18970 ;
    wire new_AGEMA_signal_18971 ;
    wire new_AGEMA_signal_18972 ;
    wire new_AGEMA_signal_18973 ;
    wire new_AGEMA_signal_18974 ;
    wire new_AGEMA_signal_18975 ;
    wire new_AGEMA_signal_18976 ;
    wire new_AGEMA_signal_18977 ;
    wire new_AGEMA_signal_18978 ;
    wire new_AGEMA_signal_18979 ;
    wire new_AGEMA_signal_18980 ;
    wire new_AGEMA_signal_18981 ;
    wire new_AGEMA_signal_18982 ;
    wire new_AGEMA_signal_18983 ;
    wire new_AGEMA_signal_18984 ;
    wire new_AGEMA_signal_18985 ;
    wire new_AGEMA_signal_18986 ;
    wire new_AGEMA_signal_18987 ;
    wire new_AGEMA_signal_18988 ;
    wire new_AGEMA_signal_18989 ;
    wire new_AGEMA_signal_18990 ;
    wire new_AGEMA_signal_18991 ;
    wire new_AGEMA_signal_18992 ;
    wire new_AGEMA_signal_18993 ;
    wire new_AGEMA_signal_18994 ;
    wire new_AGEMA_signal_18995 ;
    wire new_AGEMA_signal_18996 ;
    wire new_AGEMA_signal_18997 ;
    wire new_AGEMA_signal_18998 ;
    wire new_AGEMA_signal_18999 ;
    wire new_AGEMA_signal_19000 ;
    wire new_AGEMA_signal_19001 ;
    wire new_AGEMA_signal_19002 ;
    wire new_AGEMA_signal_19003 ;
    wire new_AGEMA_signal_19004 ;
    wire new_AGEMA_signal_19005 ;
    wire new_AGEMA_signal_19006 ;
    wire new_AGEMA_signal_19007 ;
    wire new_AGEMA_signal_19008 ;
    wire new_AGEMA_signal_19009 ;
    wire new_AGEMA_signal_19010 ;
    wire new_AGEMA_signal_19011 ;
    wire new_AGEMA_signal_19012 ;
    wire new_AGEMA_signal_19013 ;
    wire new_AGEMA_signal_19014 ;
    wire new_AGEMA_signal_19015 ;
    wire new_AGEMA_signal_19016 ;
    wire new_AGEMA_signal_19017 ;
    wire new_AGEMA_signal_19018 ;
    wire new_AGEMA_signal_19019 ;
    wire new_AGEMA_signal_19020 ;
    wire new_AGEMA_signal_19021 ;
    wire new_AGEMA_signal_19022 ;
    wire new_AGEMA_signal_19023 ;
    wire new_AGEMA_signal_19024 ;
    wire new_AGEMA_signal_19025 ;
    wire new_AGEMA_signal_19026 ;
    wire new_AGEMA_signal_19027 ;
    wire new_AGEMA_signal_19028 ;
    wire new_AGEMA_signal_19029 ;
    wire new_AGEMA_signal_19030 ;
    wire new_AGEMA_signal_19031 ;
    wire new_AGEMA_signal_19032 ;
    wire new_AGEMA_signal_19033 ;
    wire new_AGEMA_signal_19034 ;
    wire new_AGEMA_signal_19035 ;
    wire new_AGEMA_signal_19036 ;
    wire new_AGEMA_signal_19037 ;
    wire new_AGEMA_signal_19038 ;
    wire new_AGEMA_signal_19039 ;
    wire new_AGEMA_signal_19040 ;
    wire new_AGEMA_signal_19041 ;
    wire new_AGEMA_signal_19042 ;
    wire new_AGEMA_signal_19043 ;
    wire new_AGEMA_signal_19044 ;
    wire new_AGEMA_signal_19045 ;
    wire new_AGEMA_signal_19046 ;
    wire new_AGEMA_signal_19047 ;
    wire new_AGEMA_signal_19048 ;
    wire new_AGEMA_signal_19049 ;
    wire new_AGEMA_signal_19050 ;
    wire new_AGEMA_signal_19051 ;
    wire new_AGEMA_signal_19052 ;
    wire new_AGEMA_signal_19053 ;
    wire new_AGEMA_signal_19054 ;
    wire new_AGEMA_signal_19055 ;
    wire new_AGEMA_signal_19056 ;
    wire new_AGEMA_signal_19057 ;
    wire new_AGEMA_signal_19058 ;
    wire new_AGEMA_signal_19059 ;
    wire new_AGEMA_signal_19060 ;
    wire new_AGEMA_signal_19061 ;
    wire new_AGEMA_signal_19062 ;
    wire new_AGEMA_signal_19063 ;
    wire new_AGEMA_signal_19064 ;
    wire new_AGEMA_signal_19065 ;
    wire new_AGEMA_signal_19066 ;
    wire new_AGEMA_signal_19067 ;
    wire new_AGEMA_signal_19068 ;
    wire new_AGEMA_signal_19069 ;
    wire new_AGEMA_signal_19070 ;
    wire new_AGEMA_signal_19071 ;
    wire new_AGEMA_signal_19072 ;
    wire new_AGEMA_signal_19073 ;
    wire new_AGEMA_signal_19074 ;
    wire new_AGEMA_signal_19075 ;
    wire new_AGEMA_signal_19076 ;
    wire new_AGEMA_signal_19077 ;
    wire new_AGEMA_signal_19078 ;
    wire new_AGEMA_signal_19079 ;
    wire new_AGEMA_signal_19080 ;
    wire new_AGEMA_signal_19081 ;
    wire new_AGEMA_signal_19082 ;
    wire new_AGEMA_signal_19083 ;
    wire new_AGEMA_signal_19084 ;
    wire new_AGEMA_signal_19085 ;
    wire new_AGEMA_signal_19086 ;
    wire new_AGEMA_signal_19087 ;
    wire new_AGEMA_signal_19088 ;
    wire new_AGEMA_signal_19089 ;
    wire new_AGEMA_signal_19090 ;
    wire new_AGEMA_signal_19091 ;
    wire new_AGEMA_signal_19092 ;
    wire new_AGEMA_signal_19093 ;
    wire new_AGEMA_signal_19094 ;
    wire new_AGEMA_signal_19095 ;
    wire new_AGEMA_signal_19096 ;
    wire new_AGEMA_signal_19097 ;
    wire new_AGEMA_signal_19098 ;
    wire new_AGEMA_signal_19099 ;
    wire new_AGEMA_signal_19100 ;
    wire new_AGEMA_signal_19101 ;
    wire new_AGEMA_signal_19102 ;
    wire new_AGEMA_signal_19103 ;
    wire new_AGEMA_signal_19104 ;
    wire new_AGEMA_signal_19105 ;
    wire new_AGEMA_signal_19106 ;
    wire new_AGEMA_signal_19107 ;
    wire new_AGEMA_signal_19108 ;
    wire new_AGEMA_signal_19109 ;
    wire new_AGEMA_signal_19110 ;
    wire new_AGEMA_signal_19111 ;
    wire new_AGEMA_signal_19112 ;
    wire new_AGEMA_signal_19113 ;
    wire new_AGEMA_signal_19114 ;
    wire new_AGEMA_signal_19115 ;
    wire new_AGEMA_signal_19116 ;
    wire new_AGEMA_signal_19117 ;
    wire new_AGEMA_signal_19118 ;
    wire new_AGEMA_signal_19119 ;
    wire new_AGEMA_signal_19120 ;
    wire new_AGEMA_signal_19121 ;
    wire new_AGEMA_signal_19122 ;
    wire new_AGEMA_signal_19123 ;
    wire new_AGEMA_signal_19124 ;
    wire new_AGEMA_signal_19125 ;
    wire new_AGEMA_signal_19126 ;
    wire new_AGEMA_signal_19127 ;
    wire new_AGEMA_signal_19128 ;
    wire new_AGEMA_signal_19129 ;
    wire new_AGEMA_signal_19130 ;
    wire new_AGEMA_signal_19131 ;
    wire new_AGEMA_signal_19132 ;
    wire new_AGEMA_signal_19133 ;
    wire new_AGEMA_signal_19134 ;
    wire new_AGEMA_signal_19135 ;
    wire new_AGEMA_signal_19136 ;
    wire new_AGEMA_signal_19137 ;
    wire new_AGEMA_signal_19138 ;
    wire new_AGEMA_signal_19139 ;
    wire new_AGEMA_signal_19140 ;
    wire new_AGEMA_signal_19141 ;
    wire new_AGEMA_signal_19142 ;
    wire new_AGEMA_signal_19143 ;
    wire new_AGEMA_signal_19144 ;
    wire new_AGEMA_signal_19145 ;
    wire new_AGEMA_signal_19146 ;
    wire new_AGEMA_signal_19147 ;
    wire new_AGEMA_signal_19148 ;
    wire new_AGEMA_signal_19149 ;
    wire new_AGEMA_signal_19150 ;
    wire new_AGEMA_signal_19151 ;
    wire new_AGEMA_signal_19152 ;
    wire new_AGEMA_signal_19153 ;
    wire new_AGEMA_signal_19154 ;
    wire new_AGEMA_signal_19155 ;
    wire new_AGEMA_signal_19156 ;
    wire new_AGEMA_signal_19157 ;
    wire new_AGEMA_signal_19158 ;
    wire new_AGEMA_signal_19159 ;
    wire new_AGEMA_signal_19160 ;
    wire new_AGEMA_signal_19161 ;
    wire new_AGEMA_signal_19162 ;
    wire new_AGEMA_signal_19163 ;
    wire new_AGEMA_signal_19164 ;
    wire new_AGEMA_signal_19165 ;
    wire new_AGEMA_signal_19166 ;
    wire new_AGEMA_signal_19167 ;
    wire new_AGEMA_signal_19168 ;
    wire new_AGEMA_signal_19169 ;
    wire new_AGEMA_signal_19170 ;
    wire new_AGEMA_signal_19171 ;
    wire new_AGEMA_signal_19172 ;
    wire new_AGEMA_signal_19173 ;
    wire new_AGEMA_signal_19174 ;
    wire new_AGEMA_signal_19175 ;
    wire new_AGEMA_signal_19176 ;
    wire new_AGEMA_signal_19177 ;
    wire new_AGEMA_signal_19178 ;
    wire new_AGEMA_signal_19179 ;
    wire new_AGEMA_signal_19180 ;
    wire new_AGEMA_signal_19181 ;
    wire new_AGEMA_signal_19182 ;
    wire new_AGEMA_signal_19183 ;
    wire new_AGEMA_signal_19184 ;
    wire new_AGEMA_signal_19185 ;
    wire new_AGEMA_signal_19186 ;
    wire new_AGEMA_signal_19187 ;
    wire new_AGEMA_signal_19188 ;
    wire new_AGEMA_signal_19189 ;
    wire new_AGEMA_signal_19190 ;
    wire new_AGEMA_signal_19191 ;
    wire new_AGEMA_signal_19192 ;
    wire new_AGEMA_signal_19193 ;
    wire new_AGEMA_signal_19194 ;
    wire new_AGEMA_signal_19195 ;
    wire new_AGEMA_signal_19196 ;
    wire new_AGEMA_signal_19197 ;
    wire new_AGEMA_signal_19198 ;
    wire new_AGEMA_signal_19199 ;
    wire new_AGEMA_signal_19200 ;
    wire new_AGEMA_signal_19201 ;
    wire new_AGEMA_signal_19202 ;
    wire new_AGEMA_signal_19203 ;
    wire new_AGEMA_signal_19204 ;
    wire new_AGEMA_signal_19205 ;
    wire new_AGEMA_signal_19206 ;
    wire new_AGEMA_signal_19207 ;
    wire new_AGEMA_signal_19208 ;
    wire new_AGEMA_signal_19209 ;
    wire new_AGEMA_signal_19210 ;
    wire new_AGEMA_signal_19211 ;
    wire new_AGEMA_signal_19212 ;
    wire new_AGEMA_signal_19213 ;
    wire new_AGEMA_signal_19214 ;
    wire new_AGEMA_signal_19215 ;
    wire new_AGEMA_signal_19216 ;
    wire new_AGEMA_signal_19217 ;
    wire new_AGEMA_signal_19218 ;
    wire new_AGEMA_signal_19219 ;
    wire new_AGEMA_signal_19220 ;
    wire new_AGEMA_signal_19221 ;
    wire new_AGEMA_signal_19222 ;
    wire new_AGEMA_signal_19223 ;
    wire new_AGEMA_signal_19224 ;
    wire new_AGEMA_signal_19225 ;
    wire new_AGEMA_signal_19226 ;
    wire new_AGEMA_signal_19227 ;
    wire new_AGEMA_signal_19228 ;
    wire new_AGEMA_signal_19229 ;
    wire new_AGEMA_signal_19230 ;
    wire new_AGEMA_signal_19231 ;
    wire new_AGEMA_signal_19232 ;
    wire new_AGEMA_signal_19233 ;
    wire new_AGEMA_signal_19234 ;
    wire new_AGEMA_signal_19235 ;
    wire new_AGEMA_signal_19236 ;
    wire new_AGEMA_signal_19237 ;
    wire new_AGEMA_signal_19238 ;
    wire new_AGEMA_signal_19239 ;
    wire new_AGEMA_signal_19240 ;
    wire new_AGEMA_signal_19241 ;
    wire new_AGEMA_signal_19242 ;
    wire new_AGEMA_signal_19243 ;
    wire new_AGEMA_signal_19244 ;
    wire new_AGEMA_signal_19245 ;
    wire new_AGEMA_signal_19246 ;
    wire new_AGEMA_signal_19247 ;
    wire new_AGEMA_signal_19248 ;
    wire new_AGEMA_signal_19249 ;
    wire new_AGEMA_signal_19250 ;
    wire new_AGEMA_signal_19251 ;
    wire new_AGEMA_signal_19252 ;
    wire new_AGEMA_signal_19253 ;
    wire new_AGEMA_signal_19254 ;
    wire new_AGEMA_signal_19255 ;
    wire new_AGEMA_signal_19256 ;
    wire new_AGEMA_signal_19257 ;
    wire new_AGEMA_signal_19258 ;
    wire new_AGEMA_signal_19259 ;
    wire new_AGEMA_signal_19260 ;
    wire new_AGEMA_signal_19261 ;
    wire new_AGEMA_signal_19262 ;
    wire new_AGEMA_signal_19263 ;
    wire new_AGEMA_signal_19264 ;
    wire new_AGEMA_signal_19265 ;
    wire new_AGEMA_signal_19266 ;
    wire new_AGEMA_signal_19267 ;
    wire new_AGEMA_signal_19268 ;
    wire new_AGEMA_signal_19269 ;
    wire new_AGEMA_signal_19270 ;
    wire new_AGEMA_signal_19271 ;
    wire new_AGEMA_signal_19272 ;
    wire new_AGEMA_signal_19273 ;
    wire new_AGEMA_signal_19274 ;
    wire new_AGEMA_signal_19275 ;
    wire new_AGEMA_signal_19276 ;
    wire new_AGEMA_signal_19277 ;
    wire new_AGEMA_signal_19278 ;
    wire new_AGEMA_signal_19279 ;
    wire new_AGEMA_signal_19280 ;
    wire new_AGEMA_signal_19281 ;
    wire new_AGEMA_signal_19282 ;
    wire new_AGEMA_signal_19283 ;
    wire new_AGEMA_signal_19284 ;
    wire new_AGEMA_signal_19285 ;
    wire new_AGEMA_signal_19286 ;
    wire new_AGEMA_signal_19287 ;
    wire new_AGEMA_signal_19288 ;
    wire new_AGEMA_signal_19289 ;
    wire new_AGEMA_signal_19290 ;
    wire new_AGEMA_signal_19291 ;
    wire new_AGEMA_signal_19292 ;
    wire new_AGEMA_signal_19293 ;
    wire new_AGEMA_signal_19294 ;
    wire new_AGEMA_signal_19295 ;
    wire new_AGEMA_signal_19296 ;
    wire new_AGEMA_signal_19297 ;
    wire new_AGEMA_signal_19298 ;
    wire new_AGEMA_signal_19299 ;
    wire new_AGEMA_signal_19300 ;
    wire new_AGEMA_signal_19301 ;
    wire new_AGEMA_signal_19302 ;
    wire new_AGEMA_signal_19303 ;
    wire new_AGEMA_signal_19304 ;
    wire new_AGEMA_signal_19305 ;
    wire new_AGEMA_signal_19306 ;
    wire new_AGEMA_signal_19307 ;
    wire new_AGEMA_signal_19308 ;
    wire new_AGEMA_signal_19309 ;
    wire new_AGEMA_signal_19310 ;
    wire new_AGEMA_signal_19311 ;
    wire new_AGEMA_signal_19312 ;
    wire new_AGEMA_signal_19313 ;
    wire new_AGEMA_signal_19314 ;
    wire new_AGEMA_signal_19315 ;
    wire new_AGEMA_signal_19316 ;
    wire new_AGEMA_signal_19317 ;
    wire new_AGEMA_signal_19318 ;
    wire new_AGEMA_signal_19319 ;
    wire new_AGEMA_signal_19320 ;
    wire new_AGEMA_signal_19321 ;
    wire new_AGEMA_signal_19322 ;
    wire new_AGEMA_signal_19323 ;
    wire new_AGEMA_signal_19324 ;
    wire new_AGEMA_signal_19325 ;
    wire new_AGEMA_signal_19326 ;
    wire new_AGEMA_signal_19327 ;
    wire new_AGEMA_signal_19328 ;
    wire new_AGEMA_signal_19329 ;
    wire new_AGEMA_signal_19330 ;
    wire new_AGEMA_signal_19331 ;
    wire new_AGEMA_signal_19332 ;
    wire new_AGEMA_signal_19333 ;
    wire new_AGEMA_signal_19334 ;
    wire new_AGEMA_signal_19335 ;
    wire new_AGEMA_signal_19336 ;
    wire new_AGEMA_signal_19337 ;
    wire new_AGEMA_signal_19338 ;
    wire new_AGEMA_signal_19339 ;
    wire new_AGEMA_signal_19340 ;
    wire new_AGEMA_signal_19341 ;
    wire new_AGEMA_signal_19342 ;
    wire new_AGEMA_signal_19343 ;
    wire new_AGEMA_signal_19344 ;
    wire new_AGEMA_signal_19345 ;
    wire new_AGEMA_signal_19346 ;
    wire new_AGEMA_signal_19347 ;
    wire new_AGEMA_signal_19348 ;
    wire new_AGEMA_signal_19349 ;
    wire new_AGEMA_signal_19350 ;
    wire new_AGEMA_signal_19351 ;
    wire new_AGEMA_signal_19352 ;
    wire new_AGEMA_signal_19353 ;
    wire new_AGEMA_signal_19354 ;
    wire new_AGEMA_signal_19355 ;
    wire new_AGEMA_signal_19356 ;
    wire new_AGEMA_signal_19357 ;
    wire new_AGEMA_signal_19358 ;
    wire new_AGEMA_signal_19359 ;
    wire new_AGEMA_signal_19360 ;
    wire new_AGEMA_signal_19361 ;
    wire new_AGEMA_signal_19362 ;
    wire new_AGEMA_signal_19363 ;
    wire new_AGEMA_signal_19364 ;
    wire new_AGEMA_signal_19365 ;
    wire new_AGEMA_signal_19366 ;
    wire new_AGEMA_signal_19367 ;
    wire new_AGEMA_signal_19368 ;
    wire new_AGEMA_signal_19369 ;
    wire new_AGEMA_signal_19370 ;
    wire new_AGEMA_signal_19371 ;
    wire new_AGEMA_signal_19372 ;
    wire new_AGEMA_signal_19373 ;
    wire new_AGEMA_signal_19374 ;
    wire new_AGEMA_signal_19375 ;
    wire new_AGEMA_signal_19376 ;
    wire new_AGEMA_signal_19377 ;
    wire new_AGEMA_signal_19378 ;
    wire new_AGEMA_signal_19379 ;
    wire new_AGEMA_signal_19380 ;
    wire new_AGEMA_signal_19381 ;
    wire new_AGEMA_signal_19382 ;
    wire new_AGEMA_signal_19383 ;
    wire new_AGEMA_signal_19384 ;
    wire new_AGEMA_signal_19385 ;
    wire new_AGEMA_signal_19386 ;
    wire new_AGEMA_signal_19387 ;
    wire new_AGEMA_signal_19388 ;
    wire new_AGEMA_signal_19389 ;
    wire new_AGEMA_signal_19390 ;
    wire new_AGEMA_signal_19391 ;
    wire new_AGEMA_signal_19392 ;
    wire new_AGEMA_signal_19393 ;
    wire new_AGEMA_signal_19394 ;
    wire new_AGEMA_signal_19395 ;
    wire new_AGEMA_signal_19396 ;
    wire new_AGEMA_signal_19397 ;
    wire new_AGEMA_signal_19398 ;
    wire new_AGEMA_signal_19399 ;
    wire new_AGEMA_signal_19400 ;
    wire new_AGEMA_signal_19401 ;
    wire new_AGEMA_signal_19402 ;
    wire new_AGEMA_signal_19403 ;
    wire new_AGEMA_signal_19404 ;
    wire new_AGEMA_signal_19405 ;
    wire new_AGEMA_signal_19406 ;
    wire new_AGEMA_signal_19407 ;
    wire new_AGEMA_signal_19408 ;
    wire new_AGEMA_signal_19409 ;
    wire new_AGEMA_signal_19410 ;
    wire new_AGEMA_signal_19411 ;
    wire new_AGEMA_signal_19412 ;
    wire new_AGEMA_signal_19413 ;
    wire new_AGEMA_signal_19414 ;
    wire new_AGEMA_signal_19415 ;
    wire new_AGEMA_signal_19416 ;
    wire new_AGEMA_signal_19417 ;
    wire new_AGEMA_signal_19418 ;
    wire new_AGEMA_signal_19419 ;
    wire new_AGEMA_signal_19420 ;
    wire new_AGEMA_signal_19421 ;
    wire new_AGEMA_signal_19422 ;
    wire new_AGEMA_signal_19423 ;
    wire new_AGEMA_signal_19424 ;
    wire new_AGEMA_signal_19425 ;
    wire new_AGEMA_signal_19426 ;
    wire new_AGEMA_signal_19427 ;
    wire new_AGEMA_signal_19428 ;
    wire new_AGEMA_signal_19429 ;
    wire new_AGEMA_signal_19430 ;
    wire new_AGEMA_signal_19431 ;
    wire new_AGEMA_signal_19432 ;
    wire new_AGEMA_signal_19433 ;
    wire new_AGEMA_signal_19434 ;
    wire new_AGEMA_signal_19435 ;
    wire new_AGEMA_signal_19436 ;
    wire new_AGEMA_signal_19437 ;
    wire new_AGEMA_signal_19438 ;
    wire new_AGEMA_signal_19439 ;
    wire new_AGEMA_signal_19440 ;
    wire new_AGEMA_signal_19441 ;
    wire new_AGEMA_signal_19442 ;
    wire new_AGEMA_signal_19443 ;
    wire new_AGEMA_signal_19444 ;
    wire new_AGEMA_signal_19445 ;
    wire new_AGEMA_signal_19446 ;
    wire new_AGEMA_signal_19447 ;
    wire new_AGEMA_signal_19448 ;
    wire new_AGEMA_signal_19449 ;
    wire new_AGEMA_signal_19450 ;
    wire new_AGEMA_signal_19451 ;
    wire new_AGEMA_signal_19452 ;
    wire new_AGEMA_signal_19453 ;
    wire new_AGEMA_signal_19454 ;
    wire new_AGEMA_signal_19455 ;
    wire new_AGEMA_signal_19456 ;
    wire new_AGEMA_signal_19457 ;
    wire new_AGEMA_signal_19458 ;
    wire new_AGEMA_signal_19459 ;
    wire new_AGEMA_signal_19460 ;
    wire new_AGEMA_signal_19461 ;
    wire new_AGEMA_signal_19462 ;
    wire new_AGEMA_signal_19463 ;
    wire new_AGEMA_signal_19464 ;
    wire new_AGEMA_signal_19465 ;
    wire new_AGEMA_signal_19466 ;
    wire new_AGEMA_signal_19467 ;
    wire new_AGEMA_signal_19468 ;
    wire new_AGEMA_signal_19469 ;
    wire new_AGEMA_signal_19470 ;
    wire new_AGEMA_signal_19471 ;
    wire new_AGEMA_signal_19472 ;
    wire new_AGEMA_signal_19473 ;
    wire new_AGEMA_signal_19474 ;
    wire new_AGEMA_signal_19475 ;
    wire new_AGEMA_signal_19476 ;
    wire new_AGEMA_signal_19477 ;
    wire new_AGEMA_signal_19478 ;
    wire new_AGEMA_signal_19479 ;
    wire new_AGEMA_signal_19480 ;
    wire new_AGEMA_signal_19481 ;
    wire new_AGEMA_signal_19482 ;
    wire new_AGEMA_signal_19483 ;
    wire new_AGEMA_signal_19484 ;
    wire new_AGEMA_signal_19485 ;
    wire new_AGEMA_signal_19486 ;
    wire new_AGEMA_signal_19487 ;
    wire new_AGEMA_signal_19488 ;
    wire new_AGEMA_signal_19489 ;
    wire new_AGEMA_signal_19490 ;
    wire new_AGEMA_signal_19491 ;
    wire new_AGEMA_signal_19492 ;
    wire new_AGEMA_signal_19493 ;
    wire new_AGEMA_signal_19494 ;
    wire new_AGEMA_signal_19495 ;
    wire new_AGEMA_signal_19496 ;
    wire new_AGEMA_signal_19497 ;
    wire new_AGEMA_signal_19498 ;
    wire new_AGEMA_signal_19499 ;
    wire new_AGEMA_signal_19500 ;
    wire new_AGEMA_signal_19501 ;
    wire new_AGEMA_signal_19502 ;
    wire new_AGEMA_signal_19503 ;
    wire new_AGEMA_signal_19504 ;
    wire new_AGEMA_signal_19505 ;
    wire new_AGEMA_signal_19506 ;
    wire new_AGEMA_signal_19507 ;
    wire new_AGEMA_signal_19508 ;
    wire new_AGEMA_signal_19509 ;
    wire new_AGEMA_signal_19510 ;
    wire new_AGEMA_signal_19511 ;
    wire new_AGEMA_signal_19512 ;
    wire new_AGEMA_signal_19513 ;
    wire new_AGEMA_signal_19514 ;
    wire new_AGEMA_signal_19515 ;
    wire new_AGEMA_signal_19516 ;
    wire new_AGEMA_signal_19517 ;
    wire new_AGEMA_signal_19518 ;
    wire new_AGEMA_signal_19519 ;
    wire new_AGEMA_signal_19520 ;
    wire new_AGEMA_signal_19521 ;
    wire new_AGEMA_signal_19522 ;
    wire new_AGEMA_signal_19523 ;
    wire new_AGEMA_signal_19524 ;
    wire new_AGEMA_signal_19525 ;
    wire new_AGEMA_signal_19526 ;
    wire new_AGEMA_signal_19527 ;
    wire new_AGEMA_signal_19528 ;
    wire new_AGEMA_signal_19529 ;
    wire new_AGEMA_signal_19530 ;
    wire new_AGEMA_signal_19531 ;
    wire new_AGEMA_signal_19532 ;
    wire new_AGEMA_signal_19533 ;
    wire new_AGEMA_signal_19534 ;
    wire new_AGEMA_signal_19535 ;
    wire new_AGEMA_signal_19536 ;
    wire new_AGEMA_signal_19537 ;
    wire new_AGEMA_signal_19538 ;
    wire new_AGEMA_signal_19539 ;
    wire new_AGEMA_signal_19540 ;
    wire new_AGEMA_signal_19541 ;
    wire new_AGEMA_signal_19542 ;
    wire new_AGEMA_signal_19543 ;
    wire new_AGEMA_signal_19544 ;
    wire new_AGEMA_signal_19545 ;
    wire new_AGEMA_signal_19546 ;
    wire new_AGEMA_signal_19547 ;
    wire new_AGEMA_signal_19548 ;
    wire new_AGEMA_signal_19549 ;
    wire new_AGEMA_signal_19550 ;
    wire new_AGEMA_signal_19551 ;
    wire new_AGEMA_signal_19552 ;
    wire new_AGEMA_signal_19553 ;
    wire new_AGEMA_signal_19554 ;
    wire new_AGEMA_signal_19555 ;
    wire new_AGEMA_signal_19556 ;
    wire new_AGEMA_signal_19557 ;
    wire new_AGEMA_signal_19558 ;
    wire new_AGEMA_signal_19559 ;
    wire new_AGEMA_signal_19560 ;
    wire new_AGEMA_signal_19561 ;
    wire new_AGEMA_signal_19562 ;
    wire new_AGEMA_signal_19563 ;
    wire new_AGEMA_signal_19564 ;
    wire new_AGEMA_signal_19565 ;
    wire new_AGEMA_signal_19566 ;
    wire new_AGEMA_signal_19567 ;
    wire new_AGEMA_signal_19568 ;
    wire new_AGEMA_signal_19569 ;
    wire new_AGEMA_signal_19570 ;
    wire new_AGEMA_signal_19571 ;
    wire new_AGEMA_signal_19572 ;
    wire new_AGEMA_signal_19573 ;
    wire new_AGEMA_signal_19574 ;
    wire new_AGEMA_signal_19575 ;
    wire new_AGEMA_signal_19576 ;
    wire new_AGEMA_signal_19577 ;
    wire new_AGEMA_signal_19578 ;
    wire new_AGEMA_signal_19579 ;
    wire new_AGEMA_signal_19580 ;
    wire new_AGEMA_signal_19581 ;
    wire new_AGEMA_signal_19582 ;
    wire new_AGEMA_signal_19583 ;
    wire new_AGEMA_signal_19584 ;
    wire new_AGEMA_signal_19585 ;
    wire new_AGEMA_signal_19586 ;
    wire new_AGEMA_signal_19587 ;
    wire new_AGEMA_signal_19588 ;
    wire new_AGEMA_signal_19589 ;
    wire new_AGEMA_signal_19590 ;
    wire new_AGEMA_signal_19591 ;
    wire new_AGEMA_signal_19592 ;
    wire new_AGEMA_signal_19593 ;
    wire new_AGEMA_signal_19594 ;
    wire new_AGEMA_signal_19595 ;
    wire new_AGEMA_signal_19596 ;
    wire new_AGEMA_signal_19597 ;
    wire new_AGEMA_signal_19598 ;
    wire new_AGEMA_signal_19599 ;
    wire new_AGEMA_signal_19600 ;
    wire new_AGEMA_signal_19601 ;
    wire new_AGEMA_signal_19602 ;
    wire new_AGEMA_signal_19603 ;
    wire new_AGEMA_signal_19604 ;
    wire new_AGEMA_signal_19605 ;
    wire new_AGEMA_signal_19606 ;
    wire new_AGEMA_signal_19607 ;
    wire new_AGEMA_signal_19608 ;
    wire new_AGEMA_signal_19609 ;
    wire new_AGEMA_signal_19610 ;
    wire new_AGEMA_signal_19611 ;
    wire new_AGEMA_signal_19612 ;
    wire new_AGEMA_signal_19613 ;
    wire new_AGEMA_signal_19614 ;
    wire new_AGEMA_signal_19615 ;
    wire new_AGEMA_signal_19616 ;
    wire new_AGEMA_signal_19617 ;
    wire new_AGEMA_signal_19618 ;
    wire new_AGEMA_signal_19619 ;
    wire new_AGEMA_signal_19620 ;
    wire new_AGEMA_signal_19621 ;
    wire new_AGEMA_signal_19622 ;
    wire new_AGEMA_signal_19623 ;
    wire new_AGEMA_signal_19624 ;
    wire new_AGEMA_signal_19625 ;
    wire new_AGEMA_signal_19626 ;
    wire new_AGEMA_signal_19627 ;
    wire new_AGEMA_signal_19628 ;
    wire new_AGEMA_signal_19629 ;
    wire new_AGEMA_signal_19630 ;
    wire new_AGEMA_signal_19631 ;
    wire new_AGEMA_signal_19632 ;
    wire new_AGEMA_signal_19633 ;
    wire new_AGEMA_signal_19634 ;
    wire new_AGEMA_signal_19635 ;
    wire new_AGEMA_signal_19636 ;
    wire new_AGEMA_signal_19637 ;
    wire new_AGEMA_signal_19638 ;
    wire new_AGEMA_signal_19639 ;
    wire new_AGEMA_signal_19640 ;
    wire new_AGEMA_signal_19641 ;
    wire new_AGEMA_signal_19642 ;
    wire new_AGEMA_signal_19643 ;
    wire new_AGEMA_signal_19644 ;
    wire new_AGEMA_signal_19645 ;
    wire new_AGEMA_signal_19646 ;
    wire new_AGEMA_signal_19647 ;
    wire new_AGEMA_signal_19648 ;
    wire new_AGEMA_signal_19649 ;
    wire new_AGEMA_signal_19650 ;
    wire new_AGEMA_signal_19651 ;
    wire new_AGEMA_signal_19652 ;
    wire new_AGEMA_signal_19653 ;
    wire new_AGEMA_signal_19654 ;
    wire new_AGEMA_signal_19655 ;
    wire new_AGEMA_signal_19656 ;
    wire new_AGEMA_signal_19657 ;
    wire new_AGEMA_signal_19658 ;
    wire new_AGEMA_signal_19659 ;
    wire new_AGEMA_signal_19660 ;
    wire new_AGEMA_signal_19661 ;
    wire new_AGEMA_signal_19662 ;
    wire new_AGEMA_signal_19663 ;
    wire new_AGEMA_signal_19664 ;
    wire new_AGEMA_signal_19665 ;
    wire new_AGEMA_signal_19666 ;
    wire new_AGEMA_signal_19667 ;
    wire new_AGEMA_signal_19668 ;
    wire new_AGEMA_signal_19669 ;
    wire new_AGEMA_signal_19670 ;
    wire new_AGEMA_signal_19671 ;
    wire new_AGEMA_signal_19672 ;
    wire new_AGEMA_signal_19673 ;
    wire new_AGEMA_signal_19674 ;
    wire new_AGEMA_signal_19675 ;
    wire new_AGEMA_signal_19676 ;
    wire new_AGEMA_signal_19677 ;
    wire new_AGEMA_signal_19678 ;
    wire new_AGEMA_signal_19679 ;
    wire new_AGEMA_signal_19680 ;
    wire new_AGEMA_signal_19681 ;
    wire new_AGEMA_signal_19682 ;
    wire new_AGEMA_signal_19683 ;
    wire new_AGEMA_signal_19684 ;
    wire new_AGEMA_signal_19685 ;
    wire new_AGEMA_signal_19686 ;
    wire new_AGEMA_signal_19687 ;
    wire new_AGEMA_signal_19688 ;
    wire new_AGEMA_signal_19689 ;
    wire new_AGEMA_signal_19690 ;
    wire new_AGEMA_signal_19691 ;
    wire new_AGEMA_signal_19692 ;
    wire new_AGEMA_signal_19693 ;
    wire new_AGEMA_signal_19694 ;
    wire new_AGEMA_signal_19695 ;
    wire new_AGEMA_signal_19696 ;
    wire new_AGEMA_signal_19697 ;
    wire new_AGEMA_signal_19698 ;
    wire new_AGEMA_signal_19699 ;
    wire new_AGEMA_signal_19700 ;
    wire new_AGEMA_signal_19701 ;
    wire new_AGEMA_signal_19702 ;
    wire new_AGEMA_signal_19703 ;
    wire new_AGEMA_signal_19704 ;
    wire new_AGEMA_signal_19705 ;
    wire new_AGEMA_signal_19706 ;
    wire new_AGEMA_signal_19707 ;
    wire new_AGEMA_signal_19708 ;
    wire new_AGEMA_signal_19709 ;
    wire new_AGEMA_signal_19710 ;
    wire new_AGEMA_signal_19711 ;
    wire new_AGEMA_signal_19712 ;
    wire new_AGEMA_signal_19713 ;
    wire new_AGEMA_signal_19714 ;
    wire new_AGEMA_signal_19715 ;
    wire new_AGEMA_signal_19716 ;
    wire new_AGEMA_signal_19717 ;
    wire new_AGEMA_signal_19718 ;
    wire new_AGEMA_signal_19719 ;
    wire new_AGEMA_signal_19720 ;
    wire new_AGEMA_signal_19721 ;
    wire new_AGEMA_signal_19722 ;
    wire new_AGEMA_signal_19723 ;
    wire new_AGEMA_signal_19724 ;
    wire new_AGEMA_signal_19725 ;
    wire new_AGEMA_signal_19726 ;
    wire new_AGEMA_signal_19727 ;
    wire new_AGEMA_signal_19728 ;
    wire new_AGEMA_signal_19729 ;
    wire new_AGEMA_signal_19730 ;
    wire new_AGEMA_signal_19731 ;
    wire new_AGEMA_signal_19732 ;
    wire new_AGEMA_signal_19733 ;
    wire new_AGEMA_signal_19734 ;
    wire new_AGEMA_signal_19735 ;
    wire new_AGEMA_signal_19736 ;
    wire new_AGEMA_signal_19737 ;
    wire new_AGEMA_signal_19738 ;
    wire new_AGEMA_signal_19739 ;
    wire new_AGEMA_signal_19740 ;
    wire new_AGEMA_signal_19741 ;
    wire new_AGEMA_signal_19742 ;
    wire new_AGEMA_signal_19743 ;
    wire new_AGEMA_signal_19744 ;
    wire new_AGEMA_signal_19745 ;
    wire new_AGEMA_signal_19746 ;
    wire new_AGEMA_signal_19747 ;
    wire new_AGEMA_signal_19748 ;
    wire new_AGEMA_signal_19749 ;
    wire new_AGEMA_signal_19750 ;
    wire new_AGEMA_signal_19751 ;
    wire new_AGEMA_signal_19752 ;
    wire new_AGEMA_signal_19753 ;
    wire new_AGEMA_signal_19754 ;
    wire new_AGEMA_signal_19755 ;
    wire new_AGEMA_signal_19756 ;
    wire new_AGEMA_signal_19757 ;
    wire new_AGEMA_signal_19758 ;
    wire new_AGEMA_signal_19759 ;
    wire new_AGEMA_signal_19760 ;
    wire new_AGEMA_signal_19761 ;
    wire new_AGEMA_signal_19762 ;
    wire new_AGEMA_signal_19763 ;
    wire new_AGEMA_signal_19764 ;
    wire new_AGEMA_signal_19765 ;
    wire new_AGEMA_signal_19766 ;
    wire new_AGEMA_signal_19767 ;
    wire new_AGEMA_signal_19768 ;
    wire new_AGEMA_signal_19769 ;
    wire new_AGEMA_signal_19770 ;
    wire new_AGEMA_signal_19771 ;
    wire new_AGEMA_signal_19772 ;
    wire new_AGEMA_signal_19773 ;
    wire new_AGEMA_signal_19774 ;
    wire new_AGEMA_signal_19775 ;
    wire new_AGEMA_signal_19776 ;
    wire new_AGEMA_signal_19777 ;
    wire new_AGEMA_signal_19778 ;
    wire new_AGEMA_signal_19779 ;
    wire new_AGEMA_signal_19780 ;
    wire new_AGEMA_signal_19781 ;
    wire new_AGEMA_signal_19782 ;
    wire new_AGEMA_signal_19783 ;
    wire new_AGEMA_signal_19784 ;
    wire new_AGEMA_signal_19785 ;
    wire new_AGEMA_signal_19786 ;
    wire new_AGEMA_signal_19787 ;
    wire new_AGEMA_signal_19788 ;
    wire new_AGEMA_signal_19789 ;
    wire new_AGEMA_signal_19790 ;
    wire new_AGEMA_signal_19791 ;
    wire new_AGEMA_signal_19792 ;
    wire new_AGEMA_signal_19793 ;
    wire new_AGEMA_signal_19794 ;
    wire new_AGEMA_signal_19795 ;
    wire new_AGEMA_signal_19796 ;
    wire new_AGEMA_signal_19797 ;
    wire new_AGEMA_signal_19798 ;
    wire new_AGEMA_signal_19799 ;
    wire new_AGEMA_signal_19800 ;
    wire new_AGEMA_signal_19801 ;
    wire new_AGEMA_signal_19802 ;
    wire new_AGEMA_signal_19803 ;
    wire new_AGEMA_signal_19804 ;
    wire new_AGEMA_signal_19805 ;
    wire new_AGEMA_signal_19806 ;
    wire new_AGEMA_signal_19807 ;
    wire new_AGEMA_signal_19808 ;
    wire new_AGEMA_signal_19809 ;
    wire new_AGEMA_signal_19810 ;
    wire new_AGEMA_signal_19811 ;
    wire new_AGEMA_signal_19812 ;
    wire new_AGEMA_signal_19813 ;
    wire new_AGEMA_signal_19814 ;
    wire new_AGEMA_signal_19815 ;
    wire new_AGEMA_signal_19816 ;
    wire new_AGEMA_signal_19817 ;
    wire new_AGEMA_signal_19818 ;
    wire new_AGEMA_signal_19819 ;
    wire new_AGEMA_signal_19820 ;
    wire new_AGEMA_signal_19821 ;
    wire new_AGEMA_signal_19822 ;
    wire new_AGEMA_signal_19823 ;
    wire new_AGEMA_signal_19824 ;
    wire new_AGEMA_signal_19825 ;
    wire new_AGEMA_signal_19826 ;
    wire new_AGEMA_signal_19827 ;
    wire new_AGEMA_signal_19828 ;
    wire new_AGEMA_signal_19829 ;
    wire new_AGEMA_signal_19830 ;
    wire new_AGEMA_signal_19831 ;
    wire new_AGEMA_signal_19832 ;
    wire new_AGEMA_signal_19833 ;
    wire new_AGEMA_signal_19834 ;
    wire new_AGEMA_signal_19835 ;
    wire new_AGEMA_signal_19836 ;
    wire new_AGEMA_signal_19837 ;
    wire new_AGEMA_signal_19838 ;
    wire new_AGEMA_signal_19839 ;
    wire new_AGEMA_signal_19840 ;
    wire new_AGEMA_signal_19841 ;
    wire new_AGEMA_signal_19842 ;
    wire new_AGEMA_signal_19843 ;
    wire new_AGEMA_signal_19844 ;
    wire new_AGEMA_signal_19845 ;
    wire new_AGEMA_signal_19846 ;
    wire new_AGEMA_signal_19847 ;
    wire new_AGEMA_signal_19848 ;
    wire new_AGEMA_signal_19849 ;
    wire new_AGEMA_signal_19850 ;
    wire new_AGEMA_signal_19851 ;
    wire new_AGEMA_signal_19852 ;
    wire new_AGEMA_signal_19853 ;
    wire new_AGEMA_signal_19854 ;
    wire new_AGEMA_signal_19855 ;
    wire new_AGEMA_signal_19856 ;
    wire new_AGEMA_signal_19857 ;
    wire new_AGEMA_signal_19858 ;
    wire new_AGEMA_signal_19859 ;
    wire new_AGEMA_signal_19860 ;
    wire new_AGEMA_signal_19861 ;
    wire new_AGEMA_signal_19862 ;
    wire new_AGEMA_signal_19863 ;
    wire new_AGEMA_signal_19864 ;
    wire new_AGEMA_signal_19865 ;
    wire new_AGEMA_signal_19866 ;
    wire new_AGEMA_signal_19867 ;
    wire new_AGEMA_signal_19868 ;
    wire new_AGEMA_signal_19869 ;
    wire new_AGEMA_signal_19870 ;
    wire new_AGEMA_signal_19871 ;
    wire new_AGEMA_signal_19872 ;
    wire new_AGEMA_signal_19873 ;
    wire new_AGEMA_signal_19874 ;
    wire new_AGEMA_signal_19875 ;
    wire new_AGEMA_signal_19876 ;
    wire new_AGEMA_signal_19877 ;
    wire new_AGEMA_signal_19878 ;
    wire new_AGEMA_signal_19879 ;
    wire new_AGEMA_signal_19880 ;
    wire new_AGEMA_signal_19881 ;
    wire new_AGEMA_signal_19882 ;
    wire new_AGEMA_signal_19883 ;
    wire new_AGEMA_signal_19884 ;
    wire new_AGEMA_signal_19885 ;
    wire new_AGEMA_signal_19886 ;
    wire new_AGEMA_signal_19887 ;
    wire new_AGEMA_signal_19888 ;
    wire new_AGEMA_signal_19889 ;
    wire new_AGEMA_signal_19890 ;
    wire new_AGEMA_signal_19891 ;
    wire new_AGEMA_signal_19892 ;
    wire new_AGEMA_signal_19893 ;
    wire new_AGEMA_signal_19894 ;
    wire new_AGEMA_signal_19895 ;
    wire new_AGEMA_signal_19896 ;
    wire new_AGEMA_signal_19897 ;
    wire new_AGEMA_signal_19898 ;
    wire new_AGEMA_signal_19899 ;
    wire new_AGEMA_signal_19900 ;
    wire new_AGEMA_signal_19901 ;
    wire new_AGEMA_signal_19902 ;
    wire new_AGEMA_signal_19903 ;
    wire new_AGEMA_signal_19904 ;
    wire new_AGEMA_signal_19905 ;
    wire new_AGEMA_signal_19906 ;
    wire new_AGEMA_signal_19907 ;
    wire new_AGEMA_signal_19908 ;
    wire new_AGEMA_signal_19909 ;
    wire new_AGEMA_signal_19910 ;
    wire new_AGEMA_signal_19911 ;
    wire new_AGEMA_signal_19912 ;
    wire new_AGEMA_signal_19913 ;
    wire new_AGEMA_signal_19914 ;
    wire new_AGEMA_signal_19915 ;
    wire new_AGEMA_signal_19916 ;
    wire new_AGEMA_signal_19917 ;
    wire new_AGEMA_signal_19918 ;
    wire new_AGEMA_signal_19919 ;
    wire new_AGEMA_signal_19920 ;
    wire new_AGEMA_signal_19921 ;
    wire new_AGEMA_signal_19922 ;
    wire new_AGEMA_signal_19923 ;
    wire new_AGEMA_signal_19924 ;
    wire new_AGEMA_signal_19925 ;
    wire new_AGEMA_signal_19926 ;
    wire new_AGEMA_signal_19927 ;
    wire new_AGEMA_signal_19928 ;
    wire new_AGEMA_signal_19929 ;
    wire new_AGEMA_signal_19930 ;
    wire new_AGEMA_signal_19931 ;
    wire new_AGEMA_signal_19932 ;
    wire new_AGEMA_signal_19933 ;
    wire new_AGEMA_signal_19934 ;
    wire new_AGEMA_signal_19935 ;
    wire new_AGEMA_signal_19936 ;
    wire new_AGEMA_signal_19937 ;
    wire new_AGEMA_signal_19938 ;
    wire new_AGEMA_signal_19939 ;
    wire new_AGEMA_signal_19940 ;
    wire new_AGEMA_signal_19941 ;
    wire new_AGEMA_signal_19942 ;
    wire new_AGEMA_signal_19943 ;
    wire new_AGEMA_signal_19944 ;
    wire new_AGEMA_signal_19945 ;
    wire new_AGEMA_signal_19946 ;
    wire new_AGEMA_signal_19947 ;
    wire new_AGEMA_signal_19948 ;
    wire new_AGEMA_signal_19949 ;
    wire new_AGEMA_signal_19950 ;
    wire new_AGEMA_signal_19951 ;
    wire new_AGEMA_signal_19952 ;
    wire new_AGEMA_signal_19953 ;
    wire new_AGEMA_signal_19954 ;
    wire new_AGEMA_signal_19955 ;
    wire new_AGEMA_signal_19956 ;
    wire new_AGEMA_signal_19957 ;
    wire new_AGEMA_signal_19958 ;
    wire new_AGEMA_signal_19959 ;
    wire new_AGEMA_signal_19960 ;
    wire new_AGEMA_signal_19961 ;
    wire new_AGEMA_signal_19962 ;
    wire new_AGEMA_signal_19963 ;
    wire new_AGEMA_signal_19964 ;
    wire new_AGEMA_signal_19965 ;
    wire new_AGEMA_signal_19966 ;
    wire new_AGEMA_signal_19967 ;
    wire new_AGEMA_signal_19968 ;
    wire new_AGEMA_signal_19969 ;
    wire new_AGEMA_signal_19970 ;
    wire new_AGEMA_signal_19971 ;
    wire new_AGEMA_signal_19972 ;
    wire new_AGEMA_signal_19973 ;
    wire new_AGEMA_signal_19974 ;
    wire new_AGEMA_signal_19975 ;
    wire new_AGEMA_signal_19976 ;
    wire new_AGEMA_signal_19977 ;
    wire new_AGEMA_signal_19978 ;
    wire new_AGEMA_signal_19979 ;
    wire new_AGEMA_signal_19980 ;
    wire new_AGEMA_signal_19981 ;
    wire new_AGEMA_signal_19982 ;
    wire new_AGEMA_signal_19983 ;
    wire new_AGEMA_signal_19984 ;
    wire new_AGEMA_signal_19985 ;
    wire new_AGEMA_signal_19986 ;
    wire new_AGEMA_signal_19987 ;
    wire new_AGEMA_signal_19988 ;
    wire new_AGEMA_signal_19989 ;
    wire new_AGEMA_signal_19990 ;
    wire new_AGEMA_signal_19991 ;
    wire new_AGEMA_signal_19992 ;
    wire new_AGEMA_signal_19993 ;
    wire new_AGEMA_signal_19994 ;
    wire new_AGEMA_signal_19995 ;
    wire new_AGEMA_signal_19996 ;
    wire new_AGEMA_signal_19997 ;
    wire new_AGEMA_signal_19998 ;
    wire new_AGEMA_signal_19999 ;
    wire new_AGEMA_signal_20000 ;
    wire new_AGEMA_signal_20001 ;
    wire new_AGEMA_signal_20002 ;
    wire new_AGEMA_signal_20003 ;
    wire new_AGEMA_signal_20004 ;
    wire new_AGEMA_signal_20005 ;
    wire new_AGEMA_signal_20006 ;
    wire new_AGEMA_signal_20007 ;
    wire new_AGEMA_signal_20008 ;
    wire new_AGEMA_signal_20009 ;
    wire new_AGEMA_signal_20010 ;
    wire new_AGEMA_signal_20011 ;
    wire new_AGEMA_signal_20012 ;
    wire new_AGEMA_signal_20013 ;
    wire new_AGEMA_signal_20014 ;
    wire new_AGEMA_signal_20015 ;
    wire new_AGEMA_signal_20016 ;
    wire new_AGEMA_signal_20017 ;
    wire new_AGEMA_signal_20018 ;
    wire new_AGEMA_signal_20019 ;
    wire new_AGEMA_signal_20020 ;
    wire new_AGEMA_signal_20021 ;
    wire new_AGEMA_signal_20022 ;
    wire new_AGEMA_signal_20023 ;
    wire new_AGEMA_signal_20024 ;
    wire new_AGEMA_signal_20025 ;
    wire new_AGEMA_signal_20026 ;
    wire new_AGEMA_signal_20027 ;
    wire new_AGEMA_signal_20028 ;
    wire new_AGEMA_signal_20029 ;
    wire new_AGEMA_signal_20030 ;
    wire new_AGEMA_signal_20031 ;
    wire new_AGEMA_signal_20032 ;
    wire new_AGEMA_signal_20033 ;
    wire new_AGEMA_signal_20034 ;
    wire new_AGEMA_signal_20035 ;
    wire new_AGEMA_signal_20036 ;
    wire new_AGEMA_signal_20037 ;
    wire new_AGEMA_signal_20038 ;
    wire new_AGEMA_signal_20039 ;
    wire new_AGEMA_signal_20040 ;
    wire new_AGEMA_signal_20041 ;
    wire new_AGEMA_signal_20042 ;
    wire new_AGEMA_signal_20043 ;
    wire new_AGEMA_signal_20044 ;
    wire new_AGEMA_signal_20045 ;
    wire new_AGEMA_signal_20046 ;
    wire new_AGEMA_signal_20047 ;
    wire new_AGEMA_signal_20048 ;
    wire new_AGEMA_signal_20049 ;
    wire new_AGEMA_signal_20050 ;
    wire new_AGEMA_signal_20051 ;
    wire new_AGEMA_signal_20052 ;
    wire new_AGEMA_signal_20053 ;
    wire new_AGEMA_signal_20054 ;
    wire new_AGEMA_signal_20055 ;
    wire new_AGEMA_signal_20056 ;
    wire new_AGEMA_signal_20057 ;
    wire new_AGEMA_signal_20058 ;
    wire new_AGEMA_signal_20059 ;
    wire new_AGEMA_signal_20060 ;
    wire new_AGEMA_signal_20061 ;
    wire new_AGEMA_signal_20062 ;
    wire new_AGEMA_signal_20063 ;
    wire new_AGEMA_signal_20064 ;
    wire new_AGEMA_signal_20065 ;
    wire new_AGEMA_signal_20066 ;
    wire new_AGEMA_signal_20067 ;
    wire new_AGEMA_signal_20068 ;
    wire new_AGEMA_signal_20069 ;
    wire new_AGEMA_signal_20070 ;
    wire new_AGEMA_signal_20071 ;
    wire new_AGEMA_signal_20072 ;
    wire new_AGEMA_signal_20073 ;
    wire new_AGEMA_signal_20074 ;
    wire new_AGEMA_signal_20075 ;
    wire new_AGEMA_signal_20076 ;
    wire new_AGEMA_signal_20077 ;
    wire new_AGEMA_signal_20078 ;
    wire new_AGEMA_signal_20079 ;
    wire new_AGEMA_signal_20080 ;
    wire new_AGEMA_signal_20081 ;
    wire new_AGEMA_signal_20082 ;
    wire new_AGEMA_signal_20083 ;
    wire new_AGEMA_signal_20084 ;
    wire new_AGEMA_signal_20085 ;
    wire new_AGEMA_signal_20086 ;
    wire new_AGEMA_signal_20087 ;
    wire new_AGEMA_signal_20088 ;
    wire new_AGEMA_signal_20089 ;
    wire new_AGEMA_signal_20090 ;
    wire new_AGEMA_signal_20091 ;
    wire new_AGEMA_signal_20092 ;
    wire new_AGEMA_signal_20093 ;
    wire new_AGEMA_signal_20094 ;
    wire new_AGEMA_signal_20095 ;
    wire new_AGEMA_signal_20096 ;
    wire new_AGEMA_signal_20097 ;
    wire new_AGEMA_signal_20098 ;
    wire new_AGEMA_signal_20099 ;
    wire new_AGEMA_signal_20100 ;
    wire new_AGEMA_signal_20101 ;
    wire new_AGEMA_signal_20102 ;
    wire new_AGEMA_signal_20103 ;
    wire new_AGEMA_signal_20104 ;
    wire new_AGEMA_signal_20105 ;
    wire new_AGEMA_signal_20106 ;
    wire new_AGEMA_signal_20107 ;
    wire new_AGEMA_signal_20108 ;
    wire new_AGEMA_signal_20109 ;
    wire new_AGEMA_signal_20110 ;
    wire new_AGEMA_signal_20111 ;
    wire new_AGEMA_signal_20112 ;
    wire new_AGEMA_signal_20113 ;
    wire new_AGEMA_signal_20114 ;
    wire new_AGEMA_signal_20115 ;
    wire new_AGEMA_signal_20116 ;
    wire new_AGEMA_signal_20117 ;
    wire new_AGEMA_signal_20118 ;
    wire new_AGEMA_signal_20119 ;
    wire new_AGEMA_signal_20120 ;
    wire new_AGEMA_signal_20121 ;
    wire new_AGEMA_signal_20122 ;
    wire new_AGEMA_signal_20123 ;
    wire new_AGEMA_signal_20124 ;
    wire new_AGEMA_signal_20125 ;
    wire new_AGEMA_signal_20126 ;
    wire new_AGEMA_signal_20127 ;
    wire new_AGEMA_signal_20128 ;
    wire new_AGEMA_signal_20129 ;
    wire new_AGEMA_signal_20130 ;
    wire new_AGEMA_signal_20131 ;
    wire new_AGEMA_signal_20132 ;
    wire new_AGEMA_signal_20133 ;
    wire new_AGEMA_signal_20134 ;
    wire new_AGEMA_signal_20135 ;
    wire new_AGEMA_signal_20136 ;
    wire new_AGEMA_signal_20137 ;
    wire new_AGEMA_signal_20138 ;
    wire new_AGEMA_signal_20139 ;
    wire new_AGEMA_signal_20140 ;
    wire new_AGEMA_signal_20141 ;
    wire new_AGEMA_signal_20142 ;
    wire new_AGEMA_signal_20143 ;
    wire new_AGEMA_signal_20144 ;
    wire new_AGEMA_signal_20145 ;
    wire new_AGEMA_signal_20146 ;
    wire new_AGEMA_signal_20147 ;
    wire new_AGEMA_signal_20148 ;
    wire new_AGEMA_signal_20149 ;
    wire new_AGEMA_signal_20150 ;
    wire new_AGEMA_signal_20151 ;
    wire new_AGEMA_signal_20152 ;
    wire new_AGEMA_signal_20153 ;
    wire new_AGEMA_signal_20154 ;
    wire new_AGEMA_signal_20155 ;
    wire new_AGEMA_signal_20156 ;
    wire new_AGEMA_signal_20157 ;
    wire new_AGEMA_signal_20158 ;
    wire new_AGEMA_signal_20159 ;
    wire new_AGEMA_signal_20160 ;
    wire new_AGEMA_signal_20161 ;
    wire new_AGEMA_signal_20162 ;
    wire new_AGEMA_signal_20163 ;
    wire new_AGEMA_signal_20164 ;
    wire new_AGEMA_signal_20165 ;
    wire new_AGEMA_signal_20166 ;
    wire new_AGEMA_signal_20167 ;
    wire new_AGEMA_signal_20168 ;
    wire new_AGEMA_signal_20169 ;
    wire new_AGEMA_signal_20170 ;
    wire new_AGEMA_signal_20171 ;
    wire new_AGEMA_signal_20172 ;
    wire new_AGEMA_signal_20173 ;
    wire new_AGEMA_signal_20174 ;
    wire new_AGEMA_signal_20175 ;
    wire new_AGEMA_signal_20176 ;
    wire new_AGEMA_signal_20177 ;
    wire new_AGEMA_signal_20178 ;
    wire new_AGEMA_signal_20179 ;
    wire new_AGEMA_signal_20180 ;
    wire new_AGEMA_signal_20181 ;
    wire new_AGEMA_signal_20182 ;
    wire new_AGEMA_signal_20183 ;
    wire new_AGEMA_signal_20184 ;
    wire new_AGEMA_signal_20185 ;
    wire new_AGEMA_signal_20186 ;
    wire new_AGEMA_signal_20187 ;
    wire new_AGEMA_signal_20188 ;
    wire new_AGEMA_signal_20189 ;
    wire new_AGEMA_signal_20190 ;
    wire new_AGEMA_signal_20191 ;
    wire new_AGEMA_signal_20192 ;
    wire new_AGEMA_signal_20193 ;
    wire new_AGEMA_signal_20194 ;
    wire new_AGEMA_signal_20195 ;
    wire new_AGEMA_signal_20196 ;
    wire new_AGEMA_signal_20197 ;
    wire new_AGEMA_signal_20198 ;
    wire new_AGEMA_signal_20199 ;
    wire new_AGEMA_signal_20200 ;
    wire new_AGEMA_signal_20201 ;
    wire new_AGEMA_signal_20202 ;
    wire new_AGEMA_signal_20203 ;
    wire new_AGEMA_signal_20204 ;
    wire new_AGEMA_signal_20205 ;
    wire new_AGEMA_signal_20206 ;
    wire new_AGEMA_signal_20207 ;
    wire new_AGEMA_signal_20208 ;
    wire new_AGEMA_signal_20209 ;
    wire new_AGEMA_signal_20210 ;
    wire new_AGEMA_signal_20211 ;
    wire new_AGEMA_signal_20212 ;
    wire new_AGEMA_signal_20213 ;
    wire new_AGEMA_signal_20214 ;
    wire new_AGEMA_signal_20215 ;
    wire new_AGEMA_signal_20216 ;
    wire new_AGEMA_signal_20217 ;
    wire new_AGEMA_signal_20218 ;
    wire new_AGEMA_signal_20219 ;
    wire new_AGEMA_signal_20220 ;
    wire new_AGEMA_signal_20221 ;
    wire new_AGEMA_signal_20222 ;
    wire new_AGEMA_signal_20223 ;
    wire new_AGEMA_signal_20224 ;
    wire new_AGEMA_signal_20225 ;
    wire new_AGEMA_signal_20226 ;
    wire new_AGEMA_signal_20227 ;
    wire new_AGEMA_signal_20228 ;
    wire new_AGEMA_signal_20229 ;
    wire new_AGEMA_signal_20230 ;
    wire new_AGEMA_signal_20231 ;
    wire new_AGEMA_signal_20232 ;
    wire new_AGEMA_signal_20233 ;
    wire new_AGEMA_signal_20234 ;
    wire new_AGEMA_signal_20235 ;
    wire new_AGEMA_signal_20236 ;
    wire new_AGEMA_signal_20237 ;
    wire new_AGEMA_signal_20238 ;
    wire new_AGEMA_signal_20239 ;
    wire new_AGEMA_signal_20240 ;
    wire new_AGEMA_signal_20241 ;
    wire new_AGEMA_signal_20242 ;
    wire new_AGEMA_signal_20243 ;
    wire new_AGEMA_signal_20244 ;
    wire new_AGEMA_signal_20245 ;
    wire new_AGEMA_signal_20246 ;
    wire new_AGEMA_signal_20247 ;
    wire new_AGEMA_signal_20248 ;
    wire new_AGEMA_signal_20249 ;
    wire new_AGEMA_signal_20250 ;
    wire new_AGEMA_signal_20251 ;
    wire new_AGEMA_signal_20252 ;
    wire new_AGEMA_signal_20253 ;
    wire new_AGEMA_signal_20254 ;
    wire new_AGEMA_signal_20255 ;
    wire new_AGEMA_signal_20256 ;
    wire new_AGEMA_signal_20257 ;
    wire new_AGEMA_signal_20258 ;
    wire new_AGEMA_signal_20259 ;
    wire new_AGEMA_signal_20260 ;
    wire new_AGEMA_signal_20261 ;
    wire new_AGEMA_signal_20262 ;
    wire new_AGEMA_signal_20263 ;
    wire new_AGEMA_signal_20264 ;
    wire new_AGEMA_signal_20265 ;
    wire new_AGEMA_signal_20266 ;
    wire new_AGEMA_signal_20267 ;
    wire new_AGEMA_signal_20268 ;
    wire new_AGEMA_signal_20269 ;
    wire new_AGEMA_signal_20270 ;
    wire new_AGEMA_signal_20271 ;
    wire new_AGEMA_signal_20272 ;
    wire new_AGEMA_signal_20273 ;
    wire new_AGEMA_signal_20274 ;
    wire new_AGEMA_signal_20275 ;
    wire new_AGEMA_signal_20276 ;
    wire new_AGEMA_signal_20277 ;
    wire new_AGEMA_signal_20278 ;
    wire new_AGEMA_signal_20279 ;
    wire new_AGEMA_signal_20280 ;
    wire new_AGEMA_signal_20281 ;
    wire new_AGEMA_signal_20282 ;
    wire new_AGEMA_signal_20283 ;
    wire new_AGEMA_signal_20284 ;
    wire new_AGEMA_signal_20285 ;
    wire new_AGEMA_signal_20286 ;
    wire new_AGEMA_signal_20287 ;
    wire new_AGEMA_signal_20288 ;
    wire new_AGEMA_signal_20289 ;
    wire new_AGEMA_signal_20290 ;
    wire new_AGEMA_signal_20291 ;
    wire new_AGEMA_signal_20292 ;
    wire new_AGEMA_signal_20293 ;
    wire new_AGEMA_signal_20294 ;
    wire new_AGEMA_signal_20295 ;
    wire new_AGEMA_signal_20296 ;
    wire new_AGEMA_signal_20297 ;
    wire new_AGEMA_signal_20298 ;
    wire new_AGEMA_signal_20299 ;
    wire new_AGEMA_signal_20300 ;
    wire new_AGEMA_signal_20301 ;
    wire new_AGEMA_signal_20302 ;
    wire new_AGEMA_signal_20303 ;
    wire new_AGEMA_signal_20304 ;
    wire new_AGEMA_signal_20305 ;
    wire new_AGEMA_signal_20306 ;
    wire new_AGEMA_signal_20307 ;
    wire new_AGEMA_signal_20308 ;
    wire new_AGEMA_signal_20309 ;
    wire new_AGEMA_signal_20310 ;
    wire new_AGEMA_signal_20311 ;
    wire new_AGEMA_signal_20312 ;
    wire new_AGEMA_signal_20313 ;
    wire new_AGEMA_signal_20314 ;
    wire new_AGEMA_signal_20315 ;
    wire new_AGEMA_signal_20316 ;
    wire new_AGEMA_signal_20317 ;
    wire new_AGEMA_signal_20318 ;
    wire new_AGEMA_signal_20319 ;
    wire new_AGEMA_signal_20320 ;
    wire new_AGEMA_signal_20321 ;
    wire new_AGEMA_signal_20322 ;
    wire new_AGEMA_signal_20323 ;
    wire new_AGEMA_signal_20324 ;
    wire new_AGEMA_signal_20325 ;
    wire new_AGEMA_signal_20326 ;
    wire new_AGEMA_signal_20327 ;
    wire new_AGEMA_signal_20328 ;
    wire new_AGEMA_signal_20329 ;
    wire new_AGEMA_signal_20330 ;
    wire new_AGEMA_signal_20331 ;
    wire new_AGEMA_signal_20332 ;
    wire new_AGEMA_signal_20333 ;
    wire new_AGEMA_signal_20334 ;
    wire new_AGEMA_signal_20335 ;
    wire new_AGEMA_signal_20336 ;
    wire new_AGEMA_signal_20337 ;
    wire new_AGEMA_signal_20338 ;
    wire new_AGEMA_signal_20339 ;
    wire new_AGEMA_signal_20340 ;
    wire new_AGEMA_signal_20341 ;
    wire new_AGEMA_signal_20342 ;
    wire new_AGEMA_signal_20343 ;
    wire new_AGEMA_signal_20344 ;
    wire new_AGEMA_signal_20345 ;
    wire new_AGEMA_signal_20346 ;
    wire new_AGEMA_signal_20347 ;
    wire new_AGEMA_signal_20348 ;
    wire new_AGEMA_signal_20349 ;
    wire new_AGEMA_signal_20350 ;
    wire new_AGEMA_signal_20351 ;
    wire new_AGEMA_signal_20352 ;
    wire new_AGEMA_signal_20353 ;
    wire new_AGEMA_signal_20354 ;
    wire new_AGEMA_signal_20355 ;
    wire new_AGEMA_signal_20356 ;
    wire new_AGEMA_signal_20357 ;
    wire new_AGEMA_signal_20358 ;
    wire new_AGEMA_signal_20359 ;
    wire new_AGEMA_signal_20360 ;
    wire new_AGEMA_signal_20361 ;
    wire new_AGEMA_signal_20362 ;
    wire new_AGEMA_signal_20363 ;
    wire new_AGEMA_signal_20364 ;
    wire new_AGEMA_signal_20365 ;
    wire new_AGEMA_signal_20366 ;
    wire new_AGEMA_signal_20367 ;
    wire new_AGEMA_signal_20368 ;
    wire new_AGEMA_signal_20369 ;
    wire new_AGEMA_signal_20370 ;
    wire new_AGEMA_signal_20371 ;
    wire new_AGEMA_signal_20372 ;
    wire new_AGEMA_signal_20373 ;
    wire new_AGEMA_signal_20374 ;
    wire new_AGEMA_signal_20375 ;
    wire new_AGEMA_signal_20376 ;
    wire new_AGEMA_signal_20377 ;
    wire new_AGEMA_signal_20378 ;
    wire new_AGEMA_signal_20379 ;
    wire new_AGEMA_signal_20380 ;
    wire new_AGEMA_signal_20381 ;
    wire new_AGEMA_signal_20382 ;
    wire new_AGEMA_signal_20383 ;
    wire new_AGEMA_signal_20384 ;
    wire new_AGEMA_signal_20385 ;
    wire new_AGEMA_signal_20386 ;
    wire new_AGEMA_signal_20387 ;
    wire new_AGEMA_signal_20388 ;
    wire new_AGEMA_signal_20389 ;
    wire new_AGEMA_signal_20390 ;
    wire new_AGEMA_signal_20391 ;
    wire new_AGEMA_signal_20392 ;
    wire new_AGEMA_signal_20393 ;
    wire new_AGEMA_signal_20394 ;
    wire new_AGEMA_signal_20395 ;
    wire new_AGEMA_signal_20396 ;
    wire new_AGEMA_signal_20397 ;
    wire new_AGEMA_signal_20398 ;
    wire new_AGEMA_signal_20399 ;
    wire new_AGEMA_signal_20400 ;
    wire new_AGEMA_signal_20401 ;
    wire new_AGEMA_signal_20402 ;
    wire new_AGEMA_signal_20403 ;
    wire new_AGEMA_signal_20404 ;
    wire new_AGEMA_signal_20405 ;
    wire new_AGEMA_signal_20406 ;
    wire new_AGEMA_signal_20407 ;
    wire new_AGEMA_signal_20408 ;
    wire new_AGEMA_signal_20409 ;
    wire new_AGEMA_signal_20410 ;
    wire new_AGEMA_signal_20411 ;
    wire new_AGEMA_signal_20412 ;
    wire new_AGEMA_signal_20413 ;
    wire new_AGEMA_signal_20414 ;
    wire new_AGEMA_signal_20415 ;
    wire new_AGEMA_signal_20416 ;
    wire new_AGEMA_signal_20417 ;
    wire new_AGEMA_signal_20418 ;
    wire new_AGEMA_signal_20419 ;
    wire new_AGEMA_signal_20420 ;
    wire new_AGEMA_signal_20421 ;
    wire new_AGEMA_signal_20422 ;
    wire new_AGEMA_signal_20423 ;
    wire new_AGEMA_signal_20424 ;
    wire new_AGEMA_signal_20425 ;
    wire new_AGEMA_signal_20426 ;
    wire new_AGEMA_signal_20427 ;
    wire new_AGEMA_signal_20428 ;
    wire new_AGEMA_signal_20429 ;
    wire new_AGEMA_signal_20430 ;
    wire new_AGEMA_signal_20431 ;
    wire new_AGEMA_signal_20432 ;
    wire new_AGEMA_signal_20433 ;
    wire new_AGEMA_signal_20434 ;
    wire new_AGEMA_signal_20435 ;
    wire new_AGEMA_signal_20436 ;
    wire new_AGEMA_signal_20437 ;
    wire new_AGEMA_signal_20438 ;
    wire new_AGEMA_signal_20439 ;
    wire new_AGEMA_signal_20440 ;
    wire new_AGEMA_signal_20441 ;
    wire new_AGEMA_signal_20442 ;
    wire new_AGEMA_signal_20443 ;
    wire new_AGEMA_signal_20444 ;
    wire new_AGEMA_signal_20445 ;
    wire new_AGEMA_signal_20446 ;
    wire new_AGEMA_signal_20447 ;
    wire new_AGEMA_signal_20448 ;
    wire new_AGEMA_signal_20449 ;
    wire new_AGEMA_signal_20450 ;
    wire new_AGEMA_signal_20451 ;
    wire new_AGEMA_signal_20452 ;
    wire new_AGEMA_signal_20453 ;
    wire new_AGEMA_signal_20454 ;
    wire new_AGEMA_signal_20455 ;
    wire new_AGEMA_signal_20456 ;
    wire new_AGEMA_signal_20457 ;
    wire new_AGEMA_signal_20458 ;
    wire new_AGEMA_signal_20459 ;
    wire new_AGEMA_signal_20460 ;
    wire new_AGEMA_signal_20461 ;
    wire new_AGEMA_signal_20462 ;
    wire new_AGEMA_signal_20463 ;
    wire new_AGEMA_signal_20464 ;
    wire new_AGEMA_signal_20465 ;
    wire new_AGEMA_signal_20466 ;
    wire new_AGEMA_signal_20467 ;
    wire new_AGEMA_signal_20468 ;
    wire new_AGEMA_signal_20469 ;
    wire new_AGEMA_signal_20470 ;
    wire new_AGEMA_signal_20471 ;
    wire new_AGEMA_signal_20472 ;
    wire new_AGEMA_signal_20473 ;
    wire new_AGEMA_signal_20474 ;
    wire new_AGEMA_signal_20475 ;
    wire new_AGEMA_signal_20476 ;
    wire new_AGEMA_signal_20477 ;
    wire new_AGEMA_signal_20478 ;
    wire new_AGEMA_signal_20479 ;
    wire new_AGEMA_signal_20480 ;
    wire new_AGEMA_signal_20481 ;
    wire new_AGEMA_signal_20482 ;
    wire new_AGEMA_signal_20483 ;
    wire new_AGEMA_signal_20484 ;
    wire new_AGEMA_signal_20485 ;
    wire new_AGEMA_signal_20486 ;
    wire new_AGEMA_signal_20487 ;
    wire new_AGEMA_signal_20488 ;
    wire new_AGEMA_signal_20489 ;
    wire new_AGEMA_signal_20490 ;
    wire new_AGEMA_signal_20491 ;
    wire new_AGEMA_signal_20492 ;
    wire new_AGEMA_signal_20493 ;
    wire new_AGEMA_signal_20494 ;
    wire new_AGEMA_signal_20495 ;
    wire new_AGEMA_signal_20496 ;
    wire new_AGEMA_signal_20497 ;
    wire new_AGEMA_signal_20498 ;
    wire new_AGEMA_signal_20499 ;
    wire new_AGEMA_signal_20500 ;
    wire new_AGEMA_signal_20501 ;
    wire new_AGEMA_signal_20502 ;
    wire new_AGEMA_signal_20503 ;
    wire new_AGEMA_signal_20504 ;
    wire new_AGEMA_signal_20505 ;
    wire new_AGEMA_signal_20506 ;
    wire new_AGEMA_signal_20507 ;
    wire new_AGEMA_signal_20508 ;
    wire new_AGEMA_signal_20509 ;
    wire new_AGEMA_signal_20510 ;
    wire new_AGEMA_signal_20511 ;
    wire new_AGEMA_signal_20512 ;
    wire new_AGEMA_signal_20513 ;
    wire new_AGEMA_signal_20514 ;
    wire new_AGEMA_signal_20515 ;
    wire new_AGEMA_signal_20516 ;
    wire new_AGEMA_signal_20517 ;
    wire new_AGEMA_signal_20518 ;
    wire new_AGEMA_signal_20519 ;
    wire new_AGEMA_signal_20520 ;
    wire new_AGEMA_signal_20521 ;
    wire new_AGEMA_signal_20522 ;
    wire new_AGEMA_signal_20523 ;
    wire new_AGEMA_signal_20524 ;
    wire new_AGEMA_signal_20525 ;
    wire new_AGEMA_signal_20526 ;
    wire new_AGEMA_signal_20527 ;
    wire new_AGEMA_signal_20528 ;
    wire new_AGEMA_signal_20529 ;
    wire new_AGEMA_signal_20530 ;
    wire new_AGEMA_signal_20531 ;
    wire new_AGEMA_signal_20532 ;
    wire new_AGEMA_signal_20533 ;
    wire new_AGEMA_signal_20534 ;
    wire new_AGEMA_signal_20535 ;
    wire new_AGEMA_signal_20536 ;
    wire new_AGEMA_signal_20537 ;
    wire new_AGEMA_signal_20538 ;
    wire new_AGEMA_signal_20539 ;
    wire new_AGEMA_signal_20540 ;
    wire new_AGEMA_signal_20541 ;
    wire new_AGEMA_signal_20542 ;
    wire new_AGEMA_signal_20543 ;
    wire new_AGEMA_signal_20544 ;
    wire new_AGEMA_signal_20545 ;
    wire new_AGEMA_signal_20546 ;
    wire new_AGEMA_signal_20547 ;
    wire new_AGEMA_signal_20548 ;
    wire new_AGEMA_signal_20549 ;
    wire new_AGEMA_signal_20550 ;
    wire new_AGEMA_signal_20551 ;
    wire new_AGEMA_signal_20552 ;
    wire new_AGEMA_signal_20553 ;
    wire new_AGEMA_signal_20554 ;
    wire new_AGEMA_signal_20555 ;
    wire new_AGEMA_signal_20556 ;
    wire new_AGEMA_signal_20557 ;
    wire new_AGEMA_signal_20558 ;
    wire new_AGEMA_signal_20559 ;
    wire new_AGEMA_signal_20560 ;
    wire new_AGEMA_signal_20561 ;
    wire new_AGEMA_signal_20562 ;
    wire new_AGEMA_signal_20563 ;
    wire new_AGEMA_signal_20564 ;
    wire new_AGEMA_signal_20565 ;
    wire new_AGEMA_signal_20566 ;
    wire new_AGEMA_signal_20567 ;
    wire new_AGEMA_signal_20568 ;
    wire new_AGEMA_signal_20569 ;
    wire new_AGEMA_signal_20570 ;
    wire new_AGEMA_signal_20571 ;
    wire new_AGEMA_signal_20572 ;
    wire new_AGEMA_signal_20573 ;
    wire new_AGEMA_signal_20574 ;
    wire new_AGEMA_signal_20575 ;
    wire new_AGEMA_signal_20576 ;
    wire new_AGEMA_signal_20577 ;
    wire new_AGEMA_signal_20578 ;
    wire new_AGEMA_signal_20579 ;
    wire new_AGEMA_signal_20580 ;
    wire new_AGEMA_signal_20581 ;
    wire new_AGEMA_signal_20582 ;
    wire new_AGEMA_signal_20583 ;
    wire new_AGEMA_signal_20584 ;
    wire new_AGEMA_signal_20585 ;
    wire new_AGEMA_signal_20586 ;
    wire new_AGEMA_signal_20587 ;
    wire new_AGEMA_signal_20588 ;
    wire new_AGEMA_signal_20589 ;
    wire new_AGEMA_signal_20590 ;
    wire new_AGEMA_signal_20591 ;
    wire new_AGEMA_signal_20592 ;
    wire new_AGEMA_signal_20593 ;
    wire new_AGEMA_signal_20594 ;
    wire new_AGEMA_signal_20595 ;
    wire new_AGEMA_signal_20596 ;
    wire new_AGEMA_signal_20597 ;
    wire new_AGEMA_signal_20598 ;
    wire new_AGEMA_signal_20599 ;
    wire new_AGEMA_signal_20600 ;
    wire new_AGEMA_signal_20601 ;
    wire new_AGEMA_signal_20602 ;
    wire new_AGEMA_signal_20603 ;
    wire new_AGEMA_signal_20604 ;
    wire new_AGEMA_signal_20605 ;
    wire new_AGEMA_signal_20606 ;
    wire new_AGEMA_signal_20607 ;
    wire new_AGEMA_signal_20608 ;
    wire new_AGEMA_signal_20609 ;
    wire new_AGEMA_signal_20610 ;
    wire new_AGEMA_signal_20611 ;
    wire new_AGEMA_signal_20612 ;
    wire new_AGEMA_signal_20613 ;
    wire new_AGEMA_signal_20614 ;
    wire new_AGEMA_signal_20615 ;
    wire new_AGEMA_signal_20616 ;
    wire new_AGEMA_signal_20617 ;
    wire new_AGEMA_signal_20618 ;
    wire new_AGEMA_signal_20619 ;
    wire new_AGEMA_signal_20620 ;
    wire new_AGEMA_signal_20621 ;
    wire new_AGEMA_signal_20622 ;
    wire new_AGEMA_signal_20623 ;
    wire new_AGEMA_signal_20624 ;
    wire new_AGEMA_signal_20625 ;
    wire new_AGEMA_signal_20626 ;
    wire new_AGEMA_signal_20627 ;
    wire new_AGEMA_signal_20628 ;
    wire new_AGEMA_signal_20629 ;
    wire new_AGEMA_signal_20630 ;
    wire new_AGEMA_signal_20631 ;
    wire new_AGEMA_signal_20632 ;
    wire new_AGEMA_signal_20633 ;
    wire new_AGEMA_signal_20634 ;
    wire new_AGEMA_signal_20635 ;
    wire new_AGEMA_signal_20636 ;
    wire new_AGEMA_signal_20637 ;
    wire new_AGEMA_signal_20638 ;
    wire new_AGEMA_signal_20639 ;
    wire new_AGEMA_signal_20640 ;
    wire new_AGEMA_signal_20641 ;
    wire new_AGEMA_signal_20642 ;
    wire new_AGEMA_signal_20643 ;
    wire new_AGEMA_signal_20644 ;
    wire new_AGEMA_signal_20645 ;
    wire new_AGEMA_signal_20646 ;
    wire new_AGEMA_signal_20647 ;
    wire new_AGEMA_signal_20648 ;
    wire new_AGEMA_signal_20649 ;
    wire new_AGEMA_signal_20650 ;
    wire new_AGEMA_signal_20651 ;
    wire new_AGEMA_signal_20652 ;
    wire new_AGEMA_signal_20653 ;
    wire new_AGEMA_signal_20654 ;
    wire new_AGEMA_signal_20655 ;
    wire new_AGEMA_signal_20656 ;
    wire new_AGEMA_signal_20657 ;
    wire new_AGEMA_signal_20658 ;
    wire new_AGEMA_signal_20659 ;
    wire new_AGEMA_signal_20660 ;
    wire new_AGEMA_signal_20661 ;
    wire new_AGEMA_signal_20662 ;
    wire new_AGEMA_signal_20663 ;
    wire new_AGEMA_signal_20664 ;
    wire new_AGEMA_signal_20665 ;
    wire new_AGEMA_signal_20666 ;
    wire new_AGEMA_signal_20667 ;
    wire new_AGEMA_signal_20668 ;
    wire new_AGEMA_signal_20669 ;
    wire new_AGEMA_signal_20670 ;
    wire new_AGEMA_signal_20671 ;
    wire new_AGEMA_signal_20672 ;
    wire new_AGEMA_signal_20673 ;
    wire new_AGEMA_signal_20674 ;
    wire new_AGEMA_signal_20675 ;
    wire new_AGEMA_signal_20676 ;
    wire new_AGEMA_signal_20677 ;
    wire new_AGEMA_signal_20678 ;
    wire new_AGEMA_signal_20679 ;
    wire new_AGEMA_signal_20680 ;
    wire new_AGEMA_signal_20681 ;
    wire new_AGEMA_signal_20682 ;
    wire new_AGEMA_signal_20683 ;
    wire new_AGEMA_signal_20684 ;
    wire new_AGEMA_signal_20685 ;
    wire new_AGEMA_signal_20686 ;
    wire new_AGEMA_signal_20687 ;
    wire new_AGEMA_signal_20688 ;
    wire new_AGEMA_signal_20689 ;
    wire new_AGEMA_signal_20690 ;
    wire new_AGEMA_signal_20691 ;
    wire new_AGEMA_signal_20692 ;
    wire new_AGEMA_signal_20693 ;
    wire new_AGEMA_signal_20694 ;
    wire new_AGEMA_signal_20695 ;
    wire new_AGEMA_signal_20696 ;
    wire new_AGEMA_signal_20697 ;
    wire new_AGEMA_signal_20698 ;
    wire new_AGEMA_signal_20699 ;
    wire new_AGEMA_signal_20700 ;
    wire new_AGEMA_signal_20701 ;
    wire new_AGEMA_signal_20702 ;
    wire new_AGEMA_signal_20703 ;
    wire new_AGEMA_signal_20704 ;
    wire new_AGEMA_signal_20705 ;
    wire new_AGEMA_signal_20706 ;
    wire new_AGEMA_signal_20707 ;
    wire new_AGEMA_signal_20708 ;
    wire new_AGEMA_signal_20709 ;
    wire new_AGEMA_signal_20710 ;
    wire new_AGEMA_signal_20711 ;
    wire new_AGEMA_signal_20712 ;
    wire new_AGEMA_signal_20713 ;
    wire new_AGEMA_signal_20714 ;
    wire new_AGEMA_signal_20715 ;
    wire new_AGEMA_signal_20716 ;
    wire new_AGEMA_signal_20717 ;
    wire new_AGEMA_signal_20718 ;
    wire new_AGEMA_signal_20719 ;
    wire new_AGEMA_signal_20720 ;
    wire new_AGEMA_signal_20721 ;
    wire new_AGEMA_signal_20722 ;
    wire new_AGEMA_signal_20723 ;
    wire new_AGEMA_signal_20724 ;
    wire new_AGEMA_signal_20725 ;
    wire new_AGEMA_signal_20726 ;
    wire new_AGEMA_signal_20727 ;
    wire new_AGEMA_signal_20728 ;
    wire new_AGEMA_signal_20729 ;
    wire new_AGEMA_signal_20730 ;
    wire new_AGEMA_signal_20731 ;
    wire new_AGEMA_signal_20732 ;
    wire new_AGEMA_signal_20733 ;
    wire new_AGEMA_signal_20734 ;
    wire new_AGEMA_signal_20735 ;
    wire new_AGEMA_signal_20736 ;
    wire new_AGEMA_signal_20737 ;
    wire new_AGEMA_signal_20738 ;
    wire new_AGEMA_signal_20739 ;
    wire new_AGEMA_signal_20740 ;
    wire new_AGEMA_signal_20741 ;
    wire new_AGEMA_signal_20742 ;
    wire new_AGEMA_signal_20743 ;
    wire new_AGEMA_signal_20744 ;
    wire new_AGEMA_signal_20745 ;
    wire new_AGEMA_signal_20746 ;
    wire new_AGEMA_signal_20747 ;
    wire new_AGEMA_signal_20748 ;
    wire new_AGEMA_signal_20749 ;
    wire new_AGEMA_signal_20750 ;
    wire new_AGEMA_signal_20751 ;
    wire new_AGEMA_signal_20752 ;
    wire new_AGEMA_signal_20753 ;
    wire new_AGEMA_signal_20754 ;
    wire new_AGEMA_signal_20755 ;
    wire new_AGEMA_signal_20756 ;
    wire new_AGEMA_signal_20757 ;
    wire new_AGEMA_signal_20758 ;
    wire new_AGEMA_signal_20759 ;
    wire new_AGEMA_signal_20760 ;
    wire new_AGEMA_signal_20761 ;
    wire new_AGEMA_signal_20762 ;
    wire new_AGEMA_signal_20763 ;
    wire new_AGEMA_signal_20764 ;
    wire new_AGEMA_signal_20765 ;
    wire new_AGEMA_signal_20766 ;
    wire new_AGEMA_signal_20767 ;
    wire new_AGEMA_signal_20768 ;
    wire new_AGEMA_signal_20769 ;
    wire new_AGEMA_signal_20770 ;
    wire new_AGEMA_signal_20771 ;
    wire new_AGEMA_signal_20772 ;
    wire new_AGEMA_signal_20773 ;
    wire new_AGEMA_signal_20774 ;
    wire new_AGEMA_signal_20775 ;
    wire new_AGEMA_signal_20776 ;
    wire new_AGEMA_signal_20777 ;
    wire new_AGEMA_signal_20778 ;
    wire new_AGEMA_signal_20779 ;
    wire new_AGEMA_signal_20780 ;
    wire new_AGEMA_signal_20781 ;
    wire new_AGEMA_signal_20782 ;
    wire new_AGEMA_signal_20783 ;
    wire new_AGEMA_signal_20784 ;
    wire new_AGEMA_signal_20785 ;
    wire new_AGEMA_signal_20786 ;
    wire new_AGEMA_signal_20787 ;
    wire new_AGEMA_signal_20788 ;
    wire new_AGEMA_signal_20789 ;
    wire new_AGEMA_signal_20790 ;
    wire new_AGEMA_signal_20791 ;
    wire new_AGEMA_signal_20792 ;
    wire new_AGEMA_signal_20793 ;
    wire new_AGEMA_signal_20794 ;
    wire new_AGEMA_signal_20795 ;
    wire new_AGEMA_signal_20796 ;
    wire new_AGEMA_signal_20797 ;
    wire new_AGEMA_signal_20798 ;
    wire new_AGEMA_signal_20799 ;
    wire new_AGEMA_signal_20800 ;
    wire new_AGEMA_signal_20801 ;
    wire new_AGEMA_signal_20802 ;
    wire new_AGEMA_signal_20803 ;
    wire new_AGEMA_signal_20804 ;
    wire new_AGEMA_signal_20805 ;
    wire new_AGEMA_signal_20806 ;
    wire new_AGEMA_signal_20807 ;
    wire new_AGEMA_signal_20808 ;
    wire new_AGEMA_signal_20809 ;
    wire new_AGEMA_signal_20810 ;
    wire new_AGEMA_signal_20811 ;
    wire new_AGEMA_signal_20812 ;
    wire new_AGEMA_signal_20813 ;
    wire new_AGEMA_signal_20814 ;
    wire new_AGEMA_signal_20815 ;
    wire new_AGEMA_signal_20816 ;
    wire new_AGEMA_signal_20817 ;
    wire new_AGEMA_signal_20818 ;
    wire new_AGEMA_signal_20819 ;
    wire new_AGEMA_signal_20820 ;
    wire new_AGEMA_signal_20821 ;
    wire new_AGEMA_signal_20822 ;
    wire new_AGEMA_signal_20823 ;
    wire new_AGEMA_signal_20824 ;
    wire new_AGEMA_signal_20825 ;
    wire new_AGEMA_signal_20826 ;
    wire new_AGEMA_signal_20827 ;
    wire new_AGEMA_signal_20828 ;
    wire new_AGEMA_signal_20829 ;
    wire new_AGEMA_signal_20830 ;
    wire new_AGEMA_signal_20831 ;
    wire new_AGEMA_signal_20832 ;
    wire new_AGEMA_signal_20833 ;
    wire new_AGEMA_signal_20834 ;
    wire new_AGEMA_signal_20835 ;
    wire new_AGEMA_signal_20836 ;
    wire new_AGEMA_signal_20837 ;
    wire new_AGEMA_signal_20838 ;
    wire new_AGEMA_signal_20839 ;
    wire new_AGEMA_signal_20840 ;
    wire new_AGEMA_signal_20841 ;
    wire new_AGEMA_signal_20842 ;
    wire new_AGEMA_signal_20843 ;
    wire new_AGEMA_signal_20844 ;
    wire new_AGEMA_signal_20845 ;
    wire new_AGEMA_signal_20846 ;
    wire new_AGEMA_signal_20847 ;
    wire new_AGEMA_signal_20848 ;
    wire new_AGEMA_signal_20849 ;
    wire new_AGEMA_signal_20850 ;
    wire new_AGEMA_signal_20851 ;
    wire new_AGEMA_signal_20852 ;
    wire new_AGEMA_signal_20853 ;
    wire new_AGEMA_signal_20854 ;
    wire new_AGEMA_signal_20855 ;
    wire new_AGEMA_signal_20856 ;
    wire new_AGEMA_signal_20857 ;
    wire new_AGEMA_signal_20858 ;
    wire new_AGEMA_signal_20859 ;
    wire new_AGEMA_signal_20860 ;
    wire new_AGEMA_signal_20861 ;
    wire new_AGEMA_signal_20862 ;
    wire new_AGEMA_signal_20863 ;
    wire new_AGEMA_signal_20864 ;
    wire new_AGEMA_signal_20865 ;
    wire new_AGEMA_signal_20866 ;
    wire new_AGEMA_signal_20867 ;
    wire new_AGEMA_signal_20868 ;
    wire new_AGEMA_signal_20869 ;
    wire new_AGEMA_signal_20870 ;
    wire new_AGEMA_signal_20871 ;
    wire new_AGEMA_signal_20872 ;
    wire new_AGEMA_signal_20873 ;
    wire new_AGEMA_signal_20874 ;
    wire new_AGEMA_signal_20875 ;
    wire new_AGEMA_signal_20876 ;
    wire new_AGEMA_signal_20877 ;
    wire new_AGEMA_signal_20878 ;
    wire new_AGEMA_signal_20879 ;
    wire new_AGEMA_signal_20880 ;
    wire new_AGEMA_signal_20881 ;
    wire new_AGEMA_signal_20882 ;
    wire new_AGEMA_signal_20883 ;
    wire new_AGEMA_signal_20884 ;
    wire new_AGEMA_signal_20885 ;
    wire new_AGEMA_signal_20886 ;
    wire new_AGEMA_signal_20887 ;
    wire new_AGEMA_signal_20888 ;
    wire new_AGEMA_signal_20889 ;
    wire new_AGEMA_signal_20890 ;
    wire new_AGEMA_signal_20891 ;
    wire new_AGEMA_signal_20892 ;
    wire new_AGEMA_signal_20893 ;
    wire new_AGEMA_signal_20894 ;
    wire new_AGEMA_signal_20895 ;
    wire new_AGEMA_signal_20896 ;
    wire new_AGEMA_signal_20897 ;
    wire new_AGEMA_signal_20898 ;
    wire new_AGEMA_signal_20899 ;
    wire new_AGEMA_signal_20900 ;
    wire new_AGEMA_signal_20901 ;
    wire new_AGEMA_signal_20902 ;
    wire new_AGEMA_signal_20903 ;
    wire new_AGEMA_signal_20904 ;
    wire new_AGEMA_signal_20905 ;
    wire new_AGEMA_signal_20906 ;
    wire new_AGEMA_signal_20907 ;
    wire new_AGEMA_signal_20908 ;
    wire new_AGEMA_signal_20909 ;
    wire new_AGEMA_signal_20910 ;
    wire new_AGEMA_signal_20911 ;
    wire new_AGEMA_signal_20912 ;
    wire new_AGEMA_signal_20913 ;
    wire new_AGEMA_signal_20914 ;
    wire new_AGEMA_signal_20915 ;
    wire new_AGEMA_signal_20916 ;
    wire new_AGEMA_signal_20917 ;
    wire new_AGEMA_signal_20918 ;
    wire new_AGEMA_signal_20919 ;
    wire new_AGEMA_signal_20920 ;
    wire new_AGEMA_signal_20921 ;
    wire new_AGEMA_signal_20922 ;
    wire new_AGEMA_signal_20923 ;
    wire new_AGEMA_signal_20924 ;
    wire new_AGEMA_signal_20925 ;
    wire new_AGEMA_signal_20926 ;
    wire new_AGEMA_signal_20927 ;
    wire new_AGEMA_signal_20928 ;
    wire new_AGEMA_signal_20929 ;
    wire new_AGEMA_signal_20930 ;
    wire new_AGEMA_signal_20931 ;
    wire new_AGEMA_signal_20932 ;
    wire new_AGEMA_signal_20933 ;
    wire new_AGEMA_signal_20934 ;
    wire new_AGEMA_signal_20935 ;
    wire new_AGEMA_signal_20936 ;
    wire new_AGEMA_signal_20937 ;
    wire new_AGEMA_signal_20938 ;
    wire new_AGEMA_signal_20939 ;
    wire new_AGEMA_signal_20940 ;
    wire new_AGEMA_signal_20941 ;
    wire new_AGEMA_signal_20942 ;
    wire new_AGEMA_signal_20943 ;
    wire new_AGEMA_signal_20944 ;
    wire new_AGEMA_signal_20945 ;
    wire new_AGEMA_signal_20946 ;
    wire new_AGEMA_signal_20947 ;
    wire new_AGEMA_signal_20948 ;
    wire new_AGEMA_signal_20949 ;
    wire new_AGEMA_signal_20950 ;
    wire new_AGEMA_signal_20951 ;
    wire new_AGEMA_signal_20952 ;
    wire new_AGEMA_signal_20953 ;
    wire new_AGEMA_signal_20954 ;
    wire new_AGEMA_signal_20955 ;
    wire new_AGEMA_signal_20956 ;
    wire new_AGEMA_signal_20957 ;
    wire new_AGEMA_signal_20958 ;
    wire new_AGEMA_signal_20959 ;
    wire new_AGEMA_signal_20960 ;
    wire new_AGEMA_signal_20961 ;
    wire new_AGEMA_signal_20962 ;
    wire new_AGEMA_signal_20963 ;
    wire new_AGEMA_signal_20964 ;
    wire new_AGEMA_signal_20965 ;
    wire new_AGEMA_signal_20966 ;
    wire new_AGEMA_signal_20967 ;
    wire new_AGEMA_signal_20968 ;
    wire new_AGEMA_signal_20969 ;
    wire new_AGEMA_signal_20970 ;
    wire new_AGEMA_signal_20971 ;
    wire new_AGEMA_signal_20972 ;
    wire new_AGEMA_signal_20973 ;
    wire new_AGEMA_signal_20974 ;
    wire new_AGEMA_signal_20975 ;
    wire new_AGEMA_signal_20976 ;
    wire new_AGEMA_signal_20977 ;
    wire new_AGEMA_signal_20978 ;
    wire new_AGEMA_signal_20979 ;
    wire new_AGEMA_signal_20980 ;
    wire new_AGEMA_signal_20981 ;
    wire new_AGEMA_signal_20982 ;
    wire new_AGEMA_signal_20983 ;
    wire new_AGEMA_signal_20984 ;
    wire new_AGEMA_signal_20985 ;
    wire new_AGEMA_signal_20986 ;
    wire new_AGEMA_signal_20987 ;
    wire new_AGEMA_signal_20988 ;
    wire new_AGEMA_signal_20989 ;
    wire new_AGEMA_signal_20990 ;
    wire new_AGEMA_signal_20991 ;
    wire new_AGEMA_signal_20992 ;
    wire new_AGEMA_signal_20993 ;
    wire new_AGEMA_signal_20994 ;
    wire new_AGEMA_signal_20995 ;
    wire new_AGEMA_signal_20996 ;
    wire new_AGEMA_signal_20997 ;
    wire new_AGEMA_signal_20998 ;
    wire new_AGEMA_signal_20999 ;
    wire new_AGEMA_signal_21000 ;
    wire new_AGEMA_signal_21001 ;
    wire new_AGEMA_signal_21002 ;
    wire new_AGEMA_signal_21003 ;
    wire new_AGEMA_signal_21004 ;
    wire new_AGEMA_signal_21005 ;
    wire new_AGEMA_signal_21006 ;
    wire new_AGEMA_signal_21007 ;
    wire new_AGEMA_signal_21008 ;
    wire new_AGEMA_signal_21009 ;
    wire new_AGEMA_signal_21010 ;
    wire new_AGEMA_signal_21011 ;
    wire new_AGEMA_signal_21012 ;
    wire new_AGEMA_signal_21013 ;
    wire new_AGEMA_signal_21014 ;
    wire new_AGEMA_signal_21015 ;
    wire new_AGEMA_signal_21016 ;
    wire new_AGEMA_signal_21017 ;
    wire new_AGEMA_signal_21018 ;
    wire new_AGEMA_signal_21019 ;
    wire new_AGEMA_signal_21020 ;
    wire new_AGEMA_signal_21021 ;
    wire new_AGEMA_signal_21022 ;
    wire new_AGEMA_signal_21023 ;
    wire new_AGEMA_signal_21024 ;
    wire new_AGEMA_signal_21025 ;
    wire new_AGEMA_signal_21026 ;
    wire new_AGEMA_signal_21027 ;
    wire new_AGEMA_signal_21028 ;
    wire new_AGEMA_signal_21029 ;
    wire new_AGEMA_signal_21030 ;
    wire new_AGEMA_signal_21031 ;
    wire new_AGEMA_signal_21032 ;
    wire new_AGEMA_signal_21033 ;
    wire new_AGEMA_signal_21034 ;
    wire new_AGEMA_signal_21035 ;
    wire new_AGEMA_signal_21036 ;
    wire new_AGEMA_signal_21037 ;
    wire new_AGEMA_signal_21038 ;
    wire new_AGEMA_signal_21039 ;
    wire new_AGEMA_signal_21040 ;
    wire new_AGEMA_signal_21041 ;
    wire new_AGEMA_signal_21042 ;
    wire new_AGEMA_signal_21043 ;
    wire new_AGEMA_signal_21044 ;
    wire new_AGEMA_signal_21045 ;
    wire new_AGEMA_signal_21046 ;
    wire new_AGEMA_signal_21047 ;
    wire new_AGEMA_signal_21048 ;
    wire new_AGEMA_signal_21049 ;
    wire new_AGEMA_signal_21050 ;
    wire new_AGEMA_signal_21051 ;
    wire new_AGEMA_signal_21052 ;
    wire new_AGEMA_signal_21053 ;
    wire new_AGEMA_signal_21054 ;
    wire new_AGEMA_signal_21055 ;
    wire new_AGEMA_signal_21056 ;
    wire new_AGEMA_signal_21057 ;
    wire new_AGEMA_signal_21058 ;
    wire new_AGEMA_signal_21059 ;
    wire new_AGEMA_signal_21060 ;
    wire new_AGEMA_signal_21061 ;
    wire new_AGEMA_signal_21062 ;
    wire new_AGEMA_signal_21063 ;
    wire new_AGEMA_signal_21064 ;
    wire new_AGEMA_signal_21065 ;
    wire new_AGEMA_signal_21066 ;
    wire new_AGEMA_signal_21067 ;
    wire new_AGEMA_signal_21068 ;
    wire new_AGEMA_signal_21069 ;
    wire new_AGEMA_signal_21070 ;
    wire new_AGEMA_signal_21071 ;
    wire new_AGEMA_signal_21072 ;
    wire new_AGEMA_signal_21073 ;
    wire new_AGEMA_signal_21074 ;
    wire new_AGEMA_signal_21075 ;
    wire new_AGEMA_signal_21076 ;
    wire new_AGEMA_signal_21077 ;
    wire new_AGEMA_signal_21078 ;
    wire new_AGEMA_signal_21079 ;
    wire new_AGEMA_signal_21080 ;
    wire new_AGEMA_signal_21081 ;
    wire new_AGEMA_signal_21082 ;
    wire new_AGEMA_signal_21083 ;
    wire new_AGEMA_signal_21084 ;
    wire new_AGEMA_signal_21085 ;
    wire new_AGEMA_signal_21086 ;
    wire new_AGEMA_signal_21087 ;
    wire new_AGEMA_signal_21088 ;
    wire new_AGEMA_signal_21089 ;
    wire new_AGEMA_signal_21090 ;
    wire new_AGEMA_signal_21091 ;
    wire new_AGEMA_signal_21092 ;
    wire new_AGEMA_signal_21093 ;
    wire new_AGEMA_signal_21094 ;
    wire new_AGEMA_signal_21095 ;
    wire new_AGEMA_signal_21096 ;
    wire new_AGEMA_signal_21097 ;
    wire new_AGEMA_signal_21098 ;
    wire new_AGEMA_signal_21099 ;
    wire new_AGEMA_signal_21100 ;
    wire new_AGEMA_signal_21101 ;
    wire new_AGEMA_signal_21102 ;
    wire new_AGEMA_signal_21103 ;
    wire new_AGEMA_signal_21104 ;
    wire new_AGEMA_signal_21105 ;
    wire new_AGEMA_signal_21106 ;
    wire new_AGEMA_signal_21107 ;
    wire new_AGEMA_signal_21108 ;
    wire new_AGEMA_signal_21109 ;
    wire new_AGEMA_signal_21110 ;
    wire new_AGEMA_signal_21111 ;
    wire new_AGEMA_signal_21112 ;
    wire new_AGEMA_signal_21113 ;
    wire new_AGEMA_signal_21114 ;
    wire new_AGEMA_signal_21115 ;
    wire new_AGEMA_signal_21116 ;
    wire new_AGEMA_signal_21117 ;
    wire new_AGEMA_signal_21118 ;
    wire new_AGEMA_signal_21119 ;
    wire new_AGEMA_signal_21120 ;
    wire new_AGEMA_signal_21121 ;
    wire new_AGEMA_signal_21122 ;
    wire new_AGEMA_signal_21123 ;
    wire new_AGEMA_signal_21124 ;
    wire new_AGEMA_signal_21125 ;
    wire new_AGEMA_signal_21126 ;
    wire new_AGEMA_signal_21127 ;
    wire new_AGEMA_signal_21128 ;
    wire new_AGEMA_signal_21129 ;
    wire new_AGEMA_signal_21130 ;
    wire new_AGEMA_signal_21131 ;
    wire new_AGEMA_signal_21132 ;
    wire new_AGEMA_signal_21133 ;
    wire new_AGEMA_signal_21134 ;
    wire new_AGEMA_signal_21135 ;
    wire new_AGEMA_signal_21136 ;
    wire new_AGEMA_signal_21137 ;
    wire new_AGEMA_signal_21138 ;
    wire new_AGEMA_signal_21139 ;
    wire new_AGEMA_signal_21140 ;
    wire new_AGEMA_signal_21141 ;
    wire new_AGEMA_signal_21142 ;
    wire new_AGEMA_signal_21143 ;
    wire new_AGEMA_signal_21144 ;
    wire new_AGEMA_signal_21145 ;
    wire new_AGEMA_signal_21146 ;
    wire new_AGEMA_signal_21147 ;
    wire new_AGEMA_signal_21148 ;
    wire new_AGEMA_signal_21149 ;
    wire new_AGEMA_signal_21150 ;
    wire new_AGEMA_signal_21151 ;
    wire new_AGEMA_signal_21152 ;
    wire new_AGEMA_signal_21153 ;
    wire new_AGEMA_signal_21154 ;
    wire new_AGEMA_signal_21155 ;
    wire new_AGEMA_signal_21156 ;
    wire new_AGEMA_signal_21157 ;
    wire new_AGEMA_signal_21158 ;
    wire new_AGEMA_signal_21159 ;
    wire new_AGEMA_signal_21160 ;
    wire new_AGEMA_signal_21161 ;
    wire new_AGEMA_signal_21162 ;
    wire new_AGEMA_signal_21163 ;
    wire new_AGEMA_signal_21164 ;
    wire new_AGEMA_signal_21165 ;
    wire new_AGEMA_signal_21166 ;
    wire new_AGEMA_signal_21167 ;
    wire new_AGEMA_signal_21168 ;
    wire new_AGEMA_signal_21169 ;
    wire new_AGEMA_signal_21170 ;
    wire new_AGEMA_signal_21171 ;
    wire new_AGEMA_signal_21172 ;
    wire new_AGEMA_signal_21173 ;
    wire new_AGEMA_signal_21174 ;
    wire new_AGEMA_signal_21175 ;
    wire new_AGEMA_signal_21176 ;
    wire new_AGEMA_signal_21177 ;
    wire new_AGEMA_signal_21178 ;
    wire new_AGEMA_signal_21179 ;
    wire new_AGEMA_signal_21180 ;
    wire new_AGEMA_signal_21181 ;
    wire new_AGEMA_signal_21182 ;
    wire new_AGEMA_signal_21183 ;
    wire new_AGEMA_signal_21184 ;
    wire new_AGEMA_signal_21185 ;
    wire new_AGEMA_signal_21186 ;
    wire new_AGEMA_signal_21187 ;
    wire new_AGEMA_signal_21188 ;
    wire new_AGEMA_signal_21189 ;
    wire new_AGEMA_signal_21190 ;
    wire new_AGEMA_signal_21191 ;
    wire new_AGEMA_signal_21192 ;
    wire new_AGEMA_signal_21193 ;
    wire new_AGEMA_signal_21194 ;
    wire new_AGEMA_signal_21195 ;
    wire new_AGEMA_signal_21196 ;
    wire new_AGEMA_signal_21197 ;
    wire new_AGEMA_signal_21198 ;
    wire new_AGEMA_signal_21199 ;
    wire new_AGEMA_signal_21200 ;
    wire new_AGEMA_signal_21201 ;
    wire new_AGEMA_signal_21202 ;
    wire new_AGEMA_signal_21203 ;
    wire new_AGEMA_signal_21204 ;
    wire new_AGEMA_signal_21205 ;
    wire new_AGEMA_signal_21206 ;
    wire new_AGEMA_signal_21207 ;
    wire new_AGEMA_signal_21208 ;
    wire new_AGEMA_signal_21209 ;
    wire new_AGEMA_signal_21210 ;
    wire new_AGEMA_signal_21211 ;
    wire new_AGEMA_signal_21212 ;
    wire new_AGEMA_signal_21213 ;
    wire new_AGEMA_signal_21214 ;
    wire new_AGEMA_signal_21215 ;
    wire new_AGEMA_signal_21216 ;
    wire new_AGEMA_signal_21217 ;
    wire new_AGEMA_signal_21218 ;
    wire new_AGEMA_signal_21219 ;
    wire new_AGEMA_signal_21220 ;
    wire new_AGEMA_signal_21221 ;
    wire new_AGEMA_signal_21222 ;
    wire new_AGEMA_signal_21223 ;
    wire new_AGEMA_signal_21224 ;
    wire new_AGEMA_signal_21225 ;
    wire new_AGEMA_signal_21226 ;
    wire new_AGEMA_signal_21227 ;
    wire new_AGEMA_signal_21228 ;
    wire new_AGEMA_signal_21229 ;
    wire new_AGEMA_signal_21230 ;
    wire new_AGEMA_signal_21231 ;
    wire new_AGEMA_signal_21232 ;
    wire new_AGEMA_signal_21233 ;
    wire new_AGEMA_signal_21234 ;
    wire new_AGEMA_signal_21235 ;
    wire new_AGEMA_signal_21236 ;
    wire new_AGEMA_signal_21237 ;
    wire new_AGEMA_signal_21238 ;
    wire new_AGEMA_signal_21239 ;
    wire new_AGEMA_signal_21240 ;
    wire new_AGEMA_signal_21241 ;
    wire new_AGEMA_signal_21242 ;
    wire new_AGEMA_signal_21243 ;
    wire new_AGEMA_signal_21244 ;
    wire new_AGEMA_signal_21245 ;
    wire new_AGEMA_signal_21246 ;
    wire new_AGEMA_signal_21247 ;
    wire new_AGEMA_signal_21248 ;
    wire new_AGEMA_signal_21249 ;
    wire new_AGEMA_signal_21250 ;
    wire new_AGEMA_signal_21251 ;
    wire new_AGEMA_signal_21252 ;
    wire new_AGEMA_signal_21253 ;
    wire new_AGEMA_signal_21254 ;
    wire new_AGEMA_signal_21255 ;
    wire new_AGEMA_signal_21256 ;
    wire new_AGEMA_signal_21257 ;
    wire new_AGEMA_signal_21258 ;
    wire new_AGEMA_signal_21259 ;
    wire new_AGEMA_signal_21260 ;
    wire new_AGEMA_signal_21261 ;
    wire new_AGEMA_signal_21262 ;
    wire new_AGEMA_signal_21263 ;
    wire new_AGEMA_signal_21264 ;
    wire new_AGEMA_signal_21265 ;
    wire new_AGEMA_signal_21266 ;
    wire new_AGEMA_signal_21267 ;
    wire new_AGEMA_signal_21268 ;
    wire new_AGEMA_signal_21269 ;
    wire new_AGEMA_signal_21270 ;
    wire new_AGEMA_signal_21271 ;
    wire new_AGEMA_signal_21272 ;
    wire new_AGEMA_signal_21273 ;
    wire new_AGEMA_signal_21274 ;
    wire new_AGEMA_signal_21275 ;
    wire new_AGEMA_signal_21276 ;
    wire new_AGEMA_signal_21277 ;
    wire new_AGEMA_signal_21278 ;
    wire new_AGEMA_signal_21279 ;
    wire new_AGEMA_signal_21280 ;
    wire new_AGEMA_signal_21281 ;
    wire new_AGEMA_signal_21282 ;
    wire new_AGEMA_signal_21283 ;
    wire new_AGEMA_signal_21284 ;
    wire new_AGEMA_signal_21285 ;
    wire new_AGEMA_signal_21286 ;
    wire new_AGEMA_signal_21287 ;
    wire new_AGEMA_signal_21288 ;
    wire new_AGEMA_signal_21289 ;
    wire new_AGEMA_signal_21290 ;
    wire new_AGEMA_signal_21291 ;
    wire new_AGEMA_signal_21292 ;
    wire new_AGEMA_signal_21293 ;
    wire new_AGEMA_signal_21294 ;
    wire new_AGEMA_signal_21295 ;
    wire new_AGEMA_signal_21296 ;
    wire new_AGEMA_signal_21297 ;
    wire new_AGEMA_signal_21298 ;
    wire new_AGEMA_signal_21299 ;
    wire new_AGEMA_signal_21300 ;
    wire new_AGEMA_signal_21301 ;
    wire new_AGEMA_signal_21302 ;
    wire new_AGEMA_signal_21303 ;
    wire new_AGEMA_signal_21304 ;
    wire new_AGEMA_signal_21305 ;
    wire new_AGEMA_signal_21306 ;
    wire new_AGEMA_signal_21307 ;
    wire new_AGEMA_signal_21308 ;
    wire new_AGEMA_signal_21309 ;
    wire new_AGEMA_signal_21310 ;
    wire new_AGEMA_signal_21311 ;
    wire new_AGEMA_signal_21312 ;
    wire new_AGEMA_signal_21313 ;
    wire new_AGEMA_signal_21314 ;
    wire new_AGEMA_signal_21315 ;
    wire new_AGEMA_signal_21316 ;
    wire new_AGEMA_signal_21317 ;
    wire new_AGEMA_signal_21318 ;
    wire new_AGEMA_signal_21319 ;
    wire new_AGEMA_signal_21320 ;
    wire new_AGEMA_signal_21321 ;
    wire new_AGEMA_signal_21322 ;
    wire new_AGEMA_signal_21323 ;
    wire new_AGEMA_signal_21324 ;
    wire new_AGEMA_signal_21325 ;
    wire new_AGEMA_signal_21326 ;
    wire new_AGEMA_signal_21327 ;
    wire new_AGEMA_signal_21328 ;
    wire new_AGEMA_signal_21329 ;
    wire new_AGEMA_signal_21330 ;
    wire new_AGEMA_signal_21331 ;
    wire new_AGEMA_signal_21332 ;
    wire new_AGEMA_signal_21333 ;
    wire new_AGEMA_signal_21334 ;
    wire new_AGEMA_signal_21335 ;
    wire new_AGEMA_signal_21336 ;
    wire new_AGEMA_signal_21337 ;
    wire new_AGEMA_signal_21338 ;
    wire new_AGEMA_signal_21339 ;
    wire new_AGEMA_signal_21340 ;
    wire new_AGEMA_signal_21341 ;
    wire new_AGEMA_signal_21342 ;
    wire new_AGEMA_signal_21343 ;
    wire new_AGEMA_signal_21344 ;
    wire new_AGEMA_signal_21345 ;
    wire new_AGEMA_signal_21346 ;
    wire new_AGEMA_signal_21347 ;
    wire new_AGEMA_signal_21348 ;
    wire new_AGEMA_signal_21349 ;
    wire new_AGEMA_signal_21350 ;
    wire new_AGEMA_signal_21351 ;
    wire new_AGEMA_signal_21352 ;
    wire new_AGEMA_signal_21353 ;
    wire new_AGEMA_signal_21354 ;
    wire new_AGEMA_signal_21355 ;
    wire new_AGEMA_signal_21356 ;
    wire new_AGEMA_signal_21357 ;
    wire new_AGEMA_signal_21358 ;
    wire new_AGEMA_signal_21359 ;
    wire new_AGEMA_signal_21360 ;
    wire new_AGEMA_signal_21361 ;
    wire new_AGEMA_signal_21362 ;
    wire new_AGEMA_signal_21363 ;
    wire new_AGEMA_signal_21364 ;
    wire new_AGEMA_signal_21365 ;
    wire new_AGEMA_signal_21366 ;
    wire new_AGEMA_signal_21367 ;
    wire new_AGEMA_signal_21368 ;
    wire new_AGEMA_signal_21369 ;
    wire new_AGEMA_signal_21370 ;
    wire new_AGEMA_signal_21371 ;
    wire new_AGEMA_signal_21372 ;
    wire new_AGEMA_signal_21373 ;
    wire new_AGEMA_signal_21374 ;
    wire new_AGEMA_signal_21375 ;
    wire new_AGEMA_signal_21376 ;
    wire new_AGEMA_signal_21377 ;
    wire new_AGEMA_signal_21378 ;
    wire new_AGEMA_signal_21379 ;
    wire new_AGEMA_signal_21380 ;
    wire new_AGEMA_signal_21381 ;
    wire new_AGEMA_signal_21382 ;
    wire new_AGEMA_signal_21383 ;
    wire new_AGEMA_signal_21384 ;
    wire new_AGEMA_signal_21385 ;
    wire new_AGEMA_signal_21386 ;
    wire new_AGEMA_signal_21387 ;
    wire new_AGEMA_signal_21388 ;
    wire new_AGEMA_signal_21389 ;
    wire new_AGEMA_signal_21390 ;
    wire new_AGEMA_signal_21391 ;
    wire new_AGEMA_signal_21392 ;
    wire new_AGEMA_signal_21393 ;
    wire new_AGEMA_signal_21394 ;
    wire new_AGEMA_signal_21395 ;
    wire new_AGEMA_signal_21396 ;
    wire new_AGEMA_signal_21397 ;
    wire new_AGEMA_signal_21398 ;
    wire new_AGEMA_signal_21399 ;
    wire new_AGEMA_signal_21400 ;
    wire new_AGEMA_signal_21401 ;
    wire new_AGEMA_signal_21402 ;
    wire new_AGEMA_signal_21403 ;
    wire new_AGEMA_signal_21404 ;
    wire new_AGEMA_signal_21405 ;
    wire new_AGEMA_signal_21406 ;
    wire new_AGEMA_signal_21407 ;
    wire new_AGEMA_signal_21408 ;
    wire new_AGEMA_signal_21409 ;
    wire new_AGEMA_signal_21410 ;
    wire new_AGEMA_signal_21411 ;
    wire new_AGEMA_signal_21412 ;
    wire new_AGEMA_signal_21413 ;
    wire new_AGEMA_signal_21414 ;
    wire new_AGEMA_signal_21415 ;
    wire new_AGEMA_signal_21416 ;
    wire new_AGEMA_signal_21417 ;
    wire new_AGEMA_signal_21418 ;
    wire new_AGEMA_signal_21419 ;
    wire new_AGEMA_signal_21420 ;
    wire new_AGEMA_signal_21421 ;
    wire new_AGEMA_signal_21422 ;
    wire new_AGEMA_signal_21423 ;
    wire new_AGEMA_signal_21424 ;
    wire new_AGEMA_signal_21425 ;
    wire new_AGEMA_signal_21426 ;
    wire new_AGEMA_signal_21427 ;
    wire new_AGEMA_signal_21428 ;
    wire new_AGEMA_signal_21429 ;
    wire new_AGEMA_signal_21430 ;
    wire new_AGEMA_signal_21431 ;
    wire new_AGEMA_signal_21432 ;
    wire new_AGEMA_signal_21433 ;
    wire new_AGEMA_signal_21434 ;
    wire new_AGEMA_signal_21435 ;
    wire new_AGEMA_signal_21436 ;
    wire new_AGEMA_signal_21437 ;
    wire new_AGEMA_signal_21438 ;
    wire new_AGEMA_signal_21439 ;
    wire new_AGEMA_signal_21440 ;
    wire new_AGEMA_signal_21441 ;
    wire new_AGEMA_signal_21442 ;
    wire new_AGEMA_signal_21443 ;
    wire new_AGEMA_signal_21444 ;
    wire new_AGEMA_signal_21445 ;
    wire new_AGEMA_signal_21446 ;
    wire new_AGEMA_signal_21447 ;
    wire new_AGEMA_signal_21448 ;
    wire new_AGEMA_signal_21449 ;
    wire new_AGEMA_signal_21450 ;
    wire new_AGEMA_signal_21451 ;
    wire new_AGEMA_signal_21452 ;
    wire new_AGEMA_signal_21453 ;
    wire new_AGEMA_signal_21454 ;
    wire new_AGEMA_signal_21455 ;
    wire new_AGEMA_signal_21456 ;
    wire new_AGEMA_signal_21457 ;
    wire new_AGEMA_signal_21458 ;
    wire new_AGEMA_signal_21459 ;
    wire new_AGEMA_signal_21460 ;
    wire new_AGEMA_signal_21461 ;
    wire new_AGEMA_signal_21462 ;
    wire new_AGEMA_signal_21463 ;
    wire new_AGEMA_signal_21464 ;
    wire new_AGEMA_signal_21465 ;
    wire new_AGEMA_signal_21466 ;
    wire new_AGEMA_signal_21467 ;
    wire new_AGEMA_signal_21468 ;
    wire new_AGEMA_signal_21469 ;
    wire new_AGEMA_signal_21470 ;
    wire new_AGEMA_signal_21471 ;
    wire new_AGEMA_signal_21472 ;
    wire new_AGEMA_signal_21473 ;
    wire new_AGEMA_signal_21474 ;
    wire new_AGEMA_signal_21475 ;
    wire new_AGEMA_signal_21476 ;
    wire new_AGEMA_signal_21477 ;
    wire new_AGEMA_signal_21478 ;
    wire new_AGEMA_signal_21479 ;
    wire new_AGEMA_signal_21480 ;
    wire new_AGEMA_signal_21481 ;
    wire new_AGEMA_signal_21482 ;
    wire new_AGEMA_signal_21483 ;
    wire new_AGEMA_signal_21484 ;
    wire new_AGEMA_signal_21485 ;
    wire new_AGEMA_signal_21486 ;
    wire new_AGEMA_signal_21487 ;
    wire new_AGEMA_signal_21488 ;
    wire new_AGEMA_signal_21489 ;
    wire new_AGEMA_signal_21490 ;
    wire new_AGEMA_signal_21491 ;
    wire new_AGEMA_signal_21492 ;
    wire new_AGEMA_signal_21493 ;
    wire new_AGEMA_signal_21494 ;
    wire new_AGEMA_signal_21495 ;
    wire new_AGEMA_signal_21496 ;
    wire new_AGEMA_signal_21497 ;
    wire new_AGEMA_signal_21498 ;
    wire new_AGEMA_signal_21499 ;
    wire new_AGEMA_signal_21500 ;
    wire new_AGEMA_signal_21501 ;
    wire new_AGEMA_signal_21502 ;
    wire new_AGEMA_signal_21503 ;
    wire new_AGEMA_signal_21504 ;
    wire new_AGEMA_signal_21505 ;
    wire new_AGEMA_signal_21506 ;
    wire new_AGEMA_signal_21507 ;
    wire new_AGEMA_signal_21508 ;
    wire new_AGEMA_signal_21509 ;
    wire new_AGEMA_signal_21510 ;
    wire new_AGEMA_signal_21511 ;
    wire new_AGEMA_signal_21512 ;
    wire new_AGEMA_signal_21513 ;
    wire new_AGEMA_signal_21514 ;
    wire new_AGEMA_signal_21515 ;
    wire new_AGEMA_signal_21516 ;
    wire new_AGEMA_signal_21517 ;
    wire new_AGEMA_signal_21518 ;
    wire new_AGEMA_signal_21519 ;
    wire new_AGEMA_signal_21520 ;
    wire new_AGEMA_signal_21521 ;
    wire new_AGEMA_signal_21522 ;
    wire new_AGEMA_signal_21523 ;
    wire new_AGEMA_signal_21524 ;
    wire new_AGEMA_signal_21525 ;
    wire new_AGEMA_signal_21526 ;
    wire new_AGEMA_signal_21527 ;
    wire new_AGEMA_signal_21528 ;
    wire new_AGEMA_signal_21529 ;
    wire new_AGEMA_signal_21530 ;
    wire new_AGEMA_signal_21531 ;
    wire new_AGEMA_signal_21532 ;
    wire new_AGEMA_signal_21533 ;
    wire new_AGEMA_signal_21534 ;
    wire new_AGEMA_signal_21535 ;
    wire new_AGEMA_signal_21536 ;
    wire new_AGEMA_signal_21537 ;
    wire new_AGEMA_signal_21538 ;
    wire new_AGEMA_signal_21539 ;
    wire new_AGEMA_signal_21540 ;
    wire new_AGEMA_signal_21541 ;
    wire new_AGEMA_signal_21542 ;
    wire new_AGEMA_signal_21543 ;
    wire new_AGEMA_signal_21544 ;
    wire new_AGEMA_signal_21545 ;
    wire new_AGEMA_signal_21546 ;
    wire new_AGEMA_signal_21547 ;
    wire new_AGEMA_signal_21548 ;
    wire new_AGEMA_signal_21549 ;
    wire new_AGEMA_signal_21550 ;
    wire new_AGEMA_signal_21551 ;
    wire new_AGEMA_signal_21552 ;
    wire new_AGEMA_signal_21553 ;
    wire new_AGEMA_signal_21554 ;
    wire new_AGEMA_signal_21555 ;
    wire new_AGEMA_signal_21556 ;
    wire new_AGEMA_signal_21557 ;
    wire new_AGEMA_signal_21558 ;
    wire new_AGEMA_signal_21559 ;
    wire new_AGEMA_signal_21560 ;
    wire new_AGEMA_signal_21561 ;
    wire new_AGEMA_signal_21562 ;
    wire new_AGEMA_signal_21563 ;
    wire new_AGEMA_signal_21564 ;
    wire new_AGEMA_signal_21565 ;
    wire new_AGEMA_signal_21566 ;
    wire new_AGEMA_signal_21567 ;
    wire new_AGEMA_signal_21568 ;
    wire new_AGEMA_signal_21569 ;
    wire new_AGEMA_signal_21570 ;
    wire new_AGEMA_signal_21571 ;
    wire new_AGEMA_signal_21572 ;
    wire new_AGEMA_signal_21573 ;
    wire new_AGEMA_signal_21574 ;
    wire new_AGEMA_signal_21575 ;
    wire new_AGEMA_signal_21576 ;
    wire new_AGEMA_signal_21577 ;
    wire new_AGEMA_signal_21578 ;
    wire new_AGEMA_signal_21579 ;
    wire new_AGEMA_signal_21580 ;
    wire new_AGEMA_signal_21581 ;
    wire new_AGEMA_signal_21582 ;
    wire new_AGEMA_signal_21583 ;
    wire new_AGEMA_signal_21584 ;
    wire new_AGEMA_signal_21585 ;
    wire new_AGEMA_signal_21586 ;
    wire new_AGEMA_signal_21587 ;
    wire new_AGEMA_signal_21588 ;
    wire new_AGEMA_signal_21589 ;
    wire new_AGEMA_signal_21590 ;
    wire new_AGEMA_signal_21591 ;
    wire new_AGEMA_signal_21592 ;
    wire new_AGEMA_signal_21593 ;
    wire new_AGEMA_signal_21594 ;
    wire new_AGEMA_signal_21595 ;
    wire new_AGEMA_signal_21596 ;
    wire new_AGEMA_signal_21597 ;
    wire new_AGEMA_signal_21598 ;
    wire new_AGEMA_signal_21599 ;
    wire new_AGEMA_signal_21600 ;
    wire new_AGEMA_signal_21601 ;
    wire new_AGEMA_signal_21602 ;
    wire new_AGEMA_signal_21603 ;
    wire new_AGEMA_signal_21604 ;
    wire new_AGEMA_signal_21605 ;
    wire new_AGEMA_signal_21606 ;
    wire new_AGEMA_signal_21607 ;
    wire new_AGEMA_signal_21608 ;
    wire new_AGEMA_signal_21609 ;
    wire new_AGEMA_signal_21610 ;
    wire new_AGEMA_signal_21611 ;
    wire new_AGEMA_signal_21612 ;
    wire new_AGEMA_signal_21613 ;
    wire new_AGEMA_signal_21614 ;
    wire new_AGEMA_signal_21615 ;
    wire new_AGEMA_signal_21616 ;
    wire new_AGEMA_signal_21617 ;
    wire new_AGEMA_signal_21618 ;
    wire new_AGEMA_signal_21619 ;
    wire new_AGEMA_signal_21620 ;
    wire new_AGEMA_signal_21621 ;
    wire new_AGEMA_signal_21622 ;
    wire new_AGEMA_signal_21623 ;
    wire new_AGEMA_signal_21624 ;
    wire new_AGEMA_signal_21625 ;
    wire new_AGEMA_signal_21626 ;
    wire new_AGEMA_signal_21627 ;
    wire new_AGEMA_signal_21628 ;
    wire new_AGEMA_signal_21629 ;
    wire new_AGEMA_signal_21630 ;
    wire new_AGEMA_signal_21631 ;
    wire new_AGEMA_signal_21632 ;
    wire new_AGEMA_signal_21633 ;
    wire new_AGEMA_signal_21634 ;
    wire new_AGEMA_signal_21635 ;
    wire new_AGEMA_signal_21636 ;
    wire new_AGEMA_signal_21637 ;
    wire new_AGEMA_signal_21638 ;
    wire new_AGEMA_signal_21639 ;
    wire new_AGEMA_signal_21640 ;
    wire new_AGEMA_signal_21641 ;
    wire new_AGEMA_signal_21642 ;
    wire new_AGEMA_signal_21643 ;
    wire new_AGEMA_signal_21644 ;
    wire new_AGEMA_signal_21645 ;
    wire new_AGEMA_signal_21646 ;
    wire new_AGEMA_signal_21647 ;
    wire new_AGEMA_signal_21648 ;
    wire new_AGEMA_signal_21649 ;
    wire new_AGEMA_signal_21650 ;
    wire new_AGEMA_signal_21651 ;
    wire new_AGEMA_signal_21652 ;
    wire new_AGEMA_signal_21653 ;
    wire new_AGEMA_signal_21654 ;
    wire new_AGEMA_signal_21655 ;
    wire new_AGEMA_signal_21656 ;
    wire new_AGEMA_signal_21657 ;
    wire new_AGEMA_signal_21658 ;
    wire new_AGEMA_signal_21659 ;
    wire new_AGEMA_signal_21660 ;
    wire new_AGEMA_signal_21661 ;
    wire new_AGEMA_signal_21662 ;
    wire new_AGEMA_signal_21663 ;
    wire new_AGEMA_signal_21664 ;
    wire new_AGEMA_signal_21665 ;
    wire new_AGEMA_signal_21666 ;
    wire new_AGEMA_signal_21667 ;
    wire new_AGEMA_signal_21668 ;
    wire new_AGEMA_signal_21669 ;
    wire new_AGEMA_signal_21670 ;
    wire new_AGEMA_signal_21671 ;
    wire new_AGEMA_signal_21672 ;
    wire new_AGEMA_signal_21673 ;
    wire new_AGEMA_signal_21674 ;
    wire new_AGEMA_signal_21675 ;
    wire new_AGEMA_signal_21676 ;
    wire new_AGEMA_signal_21677 ;
    wire new_AGEMA_signal_21678 ;
    wire new_AGEMA_signal_21679 ;
    wire new_AGEMA_signal_21680 ;
    wire new_AGEMA_signal_21681 ;
    wire new_AGEMA_signal_21682 ;
    wire new_AGEMA_signal_21683 ;
    wire new_AGEMA_signal_21684 ;
    wire new_AGEMA_signal_21685 ;
    wire new_AGEMA_signal_21686 ;
    wire new_AGEMA_signal_21687 ;
    wire new_AGEMA_signal_21688 ;
    wire new_AGEMA_signal_21689 ;
    wire new_AGEMA_signal_21690 ;
    wire new_AGEMA_signal_21691 ;
    wire new_AGEMA_signal_21692 ;
    wire new_AGEMA_signal_21693 ;
    wire new_AGEMA_signal_21694 ;
    wire new_AGEMA_signal_21695 ;
    wire new_AGEMA_signal_21696 ;
    wire new_AGEMA_signal_21697 ;
    wire new_AGEMA_signal_21698 ;
    wire new_AGEMA_signal_21699 ;
    wire new_AGEMA_signal_21700 ;
    wire new_AGEMA_signal_21701 ;
    wire new_AGEMA_signal_21702 ;
    wire new_AGEMA_signal_21703 ;
    wire new_AGEMA_signal_21704 ;
    wire new_AGEMA_signal_21705 ;
    wire new_AGEMA_signal_21706 ;
    wire new_AGEMA_signal_21707 ;
    wire new_AGEMA_signal_21708 ;
    wire new_AGEMA_signal_21709 ;
    wire new_AGEMA_signal_21710 ;
    wire new_AGEMA_signal_21711 ;
    wire new_AGEMA_signal_21712 ;
    wire new_AGEMA_signal_21713 ;
    wire new_AGEMA_signal_21714 ;
    wire new_AGEMA_signal_21715 ;
    wire new_AGEMA_signal_21716 ;
    wire new_AGEMA_signal_21717 ;
    wire new_AGEMA_signal_21718 ;
    wire new_AGEMA_signal_21719 ;
    wire new_AGEMA_signal_21720 ;
    wire new_AGEMA_signal_21721 ;
    wire new_AGEMA_signal_21722 ;
    wire new_AGEMA_signal_21723 ;
    wire new_AGEMA_signal_21724 ;
    wire new_AGEMA_signal_21725 ;
    wire new_AGEMA_signal_21726 ;
    wire new_AGEMA_signal_21727 ;
    wire new_AGEMA_signal_21728 ;
    wire new_AGEMA_signal_21729 ;
    wire new_AGEMA_signal_21730 ;
    wire new_AGEMA_signal_21731 ;
    wire new_AGEMA_signal_21732 ;
    wire new_AGEMA_signal_21733 ;
    wire new_AGEMA_signal_21734 ;
    wire new_AGEMA_signal_21735 ;
    wire new_AGEMA_signal_21736 ;
    wire new_AGEMA_signal_21737 ;
    wire new_AGEMA_signal_21738 ;
    wire new_AGEMA_signal_21739 ;
    wire new_AGEMA_signal_21740 ;
    wire new_AGEMA_signal_21741 ;
    wire new_AGEMA_signal_21742 ;
    wire new_AGEMA_signal_21743 ;
    wire new_AGEMA_signal_21744 ;
    wire new_AGEMA_signal_21745 ;
    wire new_AGEMA_signal_21746 ;
    wire new_AGEMA_signal_21747 ;
    wire new_AGEMA_signal_21748 ;
    wire new_AGEMA_signal_21749 ;
    wire new_AGEMA_signal_21750 ;
    wire new_AGEMA_signal_21751 ;
    wire new_AGEMA_signal_21752 ;
    wire new_AGEMA_signal_21753 ;
    wire new_AGEMA_signal_21754 ;
    wire new_AGEMA_signal_21755 ;
    wire new_AGEMA_signal_21756 ;
    wire new_AGEMA_signal_21757 ;
    wire new_AGEMA_signal_21758 ;
    wire new_AGEMA_signal_21759 ;
    wire new_AGEMA_signal_21760 ;
    wire new_AGEMA_signal_21761 ;
    wire new_AGEMA_signal_21762 ;
    wire new_AGEMA_signal_21763 ;
    wire new_AGEMA_signal_21764 ;
    wire new_AGEMA_signal_21765 ;
    wire new_AGEMA_signal_21766 ;
    wire new_AGEMA_signal_21767 ;
    wire new_AGEMA_signal_21768 ;
    wire new_AGEMA_signal_21769 ;
    wire new_AGEMA_signal_21770 ;
    wire new_AGEMA_signal_21771 ;
    wire new_AGEMA_signal_21772 ;
    wire new_AGEMA_signal_21773 ;
    wire new_AGEMA_signal_21774 ;
    wire new_AGEMA_signal_21775 ;
    wire new_AGEMA_signal_21776 ;
    wire new_AGEMA_signal_21777 ;
    wire new_AGEMA_signal_21778 ;
    wire new_AGEMA_signal_21779 ;
    wire new_AGEMA_signal_21780 ;
    wire new_AGEMA_signal_21781 ;
    wire new_AGEMA_signal_21782 ;
    wire new_AGEMA_signal_21783 ;
    wire new_AGEMA_signal_21784 ;
    wire new_AGEMA_signal_21785 ;
    wire new_AGEMA_signal_21786 ;
    wire new_AGEMA_signal_21787 ;
    wire new_AGEMA_signal_21788 ;
    wire new_AGEMA_signal_21789 ;
    wire new_AGEMA_signal_21790 ;
    wire new_AGEMA_signal_21791 ;
    wire new_AGEMA_signal_21792 ;
    wire new_AGEMA_signal_21793 ;
    wire new_AGEMA_signal_21794 ;
    wire new_AGEMA_signal_21795 ;
    wire new_AGEMA_signal_21796 ;
    wire new_AGEMA_signal_21797 ;
    wire new_AGEMA_signal_21798 ;
    wire new_AGEMA_signal_21799 ;
    wire new_AGEMA_signal_21800 ;
    wire new_AGEMA_signal_21801 ;
    wire new_AGEMA_signal_21802 ;
    wire new_AGEMA_signal_21803 ;
    wire new_AGEMA_signal_21804 ;
    wire new_AGEMA_signal_21805 ;
    wire new_AGEMA_signal_21806 ;
    wire new_AGEMA_signal_21807 ;
    wire new_AGEMA_signal_21808 ;
    wire new_AGEMA_signal_21809 ;
    wire new_AGEMA_signal_21810 ;
    wire new_AGEMA_signal_21811 ;
    wire new_AGEMA_signal_21812 ;
    wire new_AGEMA_signal_21813 ;
    wire new_AGEMA_signal_21814 ;
    wire new_AGEMA_signal_21815 ;
    wire new_AGEMA_signal_21816 ;
    wire new_AGEMA_signal_21817 ;
    wire new_AGEMA_signal_21818 ;
    wire new_AGEMA_signal_21819 ;
    wire new_AGEMA_signal_21820 ;
    wire new_AGEMA_signal_21821 ;
    wire new_AGEMA_signal_21822 ;
    wire new_AGEMA_signal_21823 ;
    wire new_AGEMA_signal_21824 ;
    wire new_AGEMA_signal_21825 ;
    wire new_AGEMA_signal_21826 ;
    wire new_AGEMA_signal_21827 ;
    wire new_AGEMA_signal_21828 ;
    wire new_AGEMA_signal_21829 ;
    wire new_AGEMA_signal_21830 ;
    wire new_AGEMA_signal_21831 ;
    wire new_AGEMA_signal_21832 ;
    wire new_AGEMA_signal_21833 ;
    wire new_AGEMA_signal_21834 ;
    wire new_AGEMA_signal_21835 ;
    wire new_AGEMA_signal_21836 ;
    wire new_AGEMA_signal_21837 ;
    wire new_AGEMA_signal_21838 ;
    wire new_AGEMA_signal_21839 ;
    wire new_AGEMA_signal_21840 ;
    wire new_AGEMA_signal_21841 ;
    wire new_AGEMA_signal_21842 ;
    wire new_AGEMA_signal_21843 ;
    wire new_AGEMA_signal_21844 ;
    wire new_AGEMA_signal_21845 ;
    wire new_AGEMA_signal_21846 ;
    wire new_AGEMA_signal_21847 ;
    wire new_AGEMA_signal_21848 ;
    wire new_AGEMA_signal_21849 ;
    wire new_AGEMA_signal_21850 ;
    wire new_AGEMA_signal_21851 ;
    wire new_AGEMA_signal_21852 ;
    wire new_AGEMA_signal_21853 ;
    wire new_AGEMA_signal_21854 ;
    wire new_AGEMA_signal_21855 ;
    wire new_AGEMA_signal_21856 ;
    wire new_AGEMA_signal_21857 ;
    wire new_AGEMA_signal_21858 ;
    wire new_AGEMA_signal_21859 ;
    wire new_AGEMA_signal_21860 ;
    wire new_AGEMA_signal_21861 ;
    wire new_AGEMA_signal_21862 ;
    wire new_AGEMA_signal_21863 ;
    wire new_AGEMA_signal_21864 ;
    wire new_AGEMA_signal_21865 ;
    wire new_AGEMA_signal_21866 ;
    wire new_AGEMA_signal_21867 ;
    wire new_AGEMA_signal_21868 ;
    wire new_AGEMA_signal_21869 ;
    wire new_AGEMA_signal_21870 ;
    wire new_AGEMA_signal_21871 ;
    wire new_AGEMA_signal_21872 ;
    wire new_AGEMA_signal_21873 ;
    wire new_AGEMA_signal_21874 ;
    wire new_AGEMA_signal_21875 ;
    wire new_AGEMA_signal_21876 ;
    wire new_AGEMA_signal_21877 ;
    wire new_AGEMA_signal_21878 ;
    wire new_AGEMA_signal_21879 ;
    wire new_AGEMA_signal_21880 ;
    wire new_AGEMA_signal_21881 ;
    wire new_AGEMA_signal_21882 ;
    wire new_AGEMA_signal_21883 ;
    wire new_AGEMA_signal_21884 ;
    wire new_AGEMA_signal_21885 ;
    wire new_AGEMA_signal_21886 ;
    wire new_AGEMA_signal_21887 ;
    wire new_AGEMA_signal_21888 ;
    wire new_AGEMA_signal_21889 ;
    wire new_AGEMA_signal_21890 ;
    wire new_AGEMA_signal_21891 ;
    wire new_AGEMA_signal_21892 ;
    wire new_AGEMA_signal_21893 ;
    wire new_AGEMA_signal_21894 ;
    wire new_AGEMA_signal_21895 ;
    wire new_AGEMA_signal_21896 ;
    wire new_AGEMA_signal_21897 ;
    wire new_AGEMA_signal_21898 ;
    wire new_AGEMA_signal_21899 ;
    wire new_AGEMA_signal_21900 ;
    wire new_AGEMA_signal_21901 ;
    wire new_AGEMA_signal_21902 ;
    wire new_AGEMA_signal_21903 ;
    wire new_AGEMA_signal_21904 ;
    wire new_AGEMA_signal_21905 ;
    wire new_AGEMA_signal_21906 ;
    wire new_AGEMA_signal_21907 ;
    wire new_AGEMA_signal_21908 ;
    wire new_AGEMA_signal_21909 ;
    wire new_AGEMA_signal_21910 ;
    wire new_AGEMA_signal_21911 ;
    wire new_AGEMA_signal_21912 ;
    wire new_AGEMA_signal_21913 ;
    wire new_AGEMA_signal_21914 ;
    wire new_AGEMA_signal_21915 ;
    wire new_AGEMA_signal_21916 ;
    wire new_AGEMA_signal_21917 ;
    wire new_AGEMA_signal_21918 ;
    wire new_AGEMA_signal_21919 ;
    wire new_AGEMA_signal_21920 ;
    wire new_AGEMA_signal_21921 ;
    wire new_AGEMA_signal_21922 ;
    wire new_AGEMA_signal_21923 ;
    wire new_AGEMA_signal_21924 ;
    wire new_AGEMA_signal_21925 ;
    wire new_AGEMA_signal_21926 ;
    wire new_AGEMA_signal_21927 ;
    wire new_AGEMA_signal_21928 ;
    wire new_AGEMA_signal_21929 ;
    wire new_AGEMA_signal_21930 ;
    wire new_AGEMA_signal_21931 ;
    wire new_AGEMA_signal_21932 ;
    wire new_AGEMA_signal_21933 ;
    wire new_AGEMA_signal_21934 ;
    wire new_AGEMA_signal_21935 ;
    wire new_AGEMA_signal_21936 ;
    wire new_AGEMA_signal_21937 ;
    wire new_AGEMA_signal_21938 ;
    wire new_AGEMA_signal_21939 ;
    wire new_AGEMA_signal_21940 ;
    wire new_AGEMA_signal_21941 ;
    wire new_AGEMA_signal_21942 ;
    wire new_AGEMA_signal_21943 ;
    wire new_AGEMA_signal_21944 ;
    wire new_AGEMA_signal_21945 ;
    wire new_AGEMA_signal_21946 ;
    wire new_AGEMA_signal_21947 ;
    wire new_AGEMA_signal_21948 ;
    wire new_AGEMA_signal_21949 ;
    wire new_AGEMA_signal_21950 ;
    wire new_AGEMA_signal_21951 ;
    wire new_AGEMA_signal_21952 ;
    wire new_AGEMA_signal_21953 ;
    wire new_AGEMA_signal_21954 ;
    wire new_AGEMA_signal_21955 ;
    wire new_AGEMA_signal_21956 ;
    wire new_AGEMA_signal_21957 ;
    wire new_AGEMA_signal_21958 ;
    wire new_AGEMA_signal_21959 ;
    wire new_AGEMA_signal_21960 ;
    wire new_AGEMA_signal_21961 ;
    wire new_AGEMA_signal_21962 ;
    wire new_AGEMA_signal_21963 ;
    wire new_AGEMA_signal_21964 ;
    wire new_AGEMA_signal_21965 ;
    wire new_AGEMA_signal_21966 ;
    wire new_AGEMA_signal_21967 ;
    wire new_AGEMA_signal_21968 ;
    wire new_AGEMA_signal_21969 ;
    wire new_AGEMA_signal_21970 ;
    wire new_AGEMA_signal_21971 ;
    wire new_AGEMA_signal_21972 ;
    wire new_AGEMA_signal_21973 ;
    wire new_AGEMA_signal_21974 ;
    wire new_AGEMA_signal_21975 ;
    wire new_AGEMA_signal_21976 ;
    wire new_AGEMA_signal_21977 ;
    wire new_AGEMA_signal_21978 ;
    wire new_AGEMA_signal_21979 ;
    wire new_AGEMA_signal_21980 ;
    wire new_AGEMA_signal_21981 ;
    wire new_AGEMA_signal_21982 ;
    wire new_AGEMA_signal_21983 ;
    wire new_AGEMA_signal_21984 ;
    wire new_AGEMA_signal_21985 ;
    wire new_AGEMA_signal_21986 ;
    wire new_AGEMA_signal_21987 ;
    wire new_AGEMA_signal_21988 ;
    wire new_AGEMA_signal_21989 ;
    wire new_AGEMA_signal_21990 ;
    wire new_AGEMA_signal_21991 ;
    wire new_AGEMA_signal_21992 ;
    wire new_AGEMA_signal_21993 ;
    wire new_AGEMA_signal_21994 ;
    wire new_AGEMA_signal_21995 ;
    wire new_AGEMA_signal_21996 ;
    wire new_AGEMA_signal_21997 ;
    wire new_AGEMA_signal_21998 ;
    wire new_AGEMA_signal_21999 ;
    wire new_AGEMA_signal_22000 ;
    wire new_AGEMA_signal_22001 ;
    wire new_AGEMA_signal_22002 ;
    wire new_AGEMA_signal_22003 ;
    wire new_AGEMA_signal_22004 ;
    wire new_AGEMA_signal_22005 ;
    wire new_AGEMA_signal_22006 ;
    wire new_AGEMA_signal_22007 ;
    wire new_AGEMA_signal_22008 ;
    wire new_AGEMA_signal_22009 ;
    wire new_AGEMA_signal_22010 ;
    wire new_AGEMA_signal_22011 ;
    wire new_AGEMA_signal_22012 ;
    wire new_AGEMA_signal_22013 ;
    wire new_AGEMA_signal_22014 ;
    wire new_AGEMA_signal_22015 ;
    wire new_AGEMA_signal_22016 ;
    wire new_AGEMA_signal_22017 ;
    wire new_AGEMA_signal_22018 ;
    wire new_AGEMA_signal_22019 ;
    wire new_AGEMA_signal_22020 ;
    wire new_AGEMA_signal_22021 ;
    wire new_AGEMA_signal_22022 ;
    wire new_AGEMA_signal_22023 ;
    wire new_AGEMA_signal_22024 ;
    wire new_AGEMA_signal_22025 ;
    wire new_AGEMA_signal_22026 ;
    wire new_AGEMA_signal_22027 ;
    wire new_AGEMA_signal_22028 ;
    wire new_AGEMA_signal_22029 ;
    wire new_AGEMA_signal_22030 ;
    wire new_AGEMA_signal_22031 ;
    wire new_AGEMA_signal_22032 ;
    wire new_AGEMA_signal_22033 ;
    wire new_AGEMA_signal_22034 ;
    wire new_AGEMA_signal_22035 ;
    wire new_AGEMA_signal_22036 ;
    wire new_AGEMA_signal_22037 ;
    wire new_AGEMA_signal_22038 ;
    wire new_AGEMA_signal_22039 ;
    wire new_AGEMA_signal_22040 ;
    wire new_AGEMA_signal_22041 ;
    wire new_AGEMA_signal_22042 ;
    wire new_AGEMA_signal_22043 ;
    wire new_AGEMA_signal_22044 ;
    wire new_AGEMA_signal_22045 ;
    wire new_AGEMA_signal_22046 ;
    wire new_AGEMA_signal_22047 ;
    wire new_AGEMA_signal_22048 ;
    wire new_AGEMA_signal_22049 ;
    wire new_AGEMA_signal_22050 ;
    wire new_AGEMA_signal_22051 ;
    wire new_AGEMA_signal_22052 ;
    wire new_AGEMA_signal_22053 ;
    wire new_AGEMA_signal_22054 ;
    wire new_AGEMA_signal_22055 ;
    wire new_AGEMA_signal_22056 ;
    wire new_AGEMA_signal_22057 ;
    wire new_AGEMA_signal_22058 ;
    wire new_AGEMA_signal_22059 ;
    wire new_AGEMA_signal_22060 ;
    wire new_AGEMA_signal_22061 ;
    wire new_AGEMA_signal_22062 ;
    wire new_AGEMA_signal_22063 ;
    wire new_AGEMA_signal_22064 ;
    wire new_AGEMA_signal_22065 ;
    wire new_AGEMA_signal_22066 ;
    wire new_AGEMA_signal_22067 ;
    wire new_AGEMA_signal_22068 ;
    wire new_AGEMA_signal_22069 ;
    wire new_AGEMA_signal_22070 ;
    wire new_AGEMA_signal_22071 ;
    wire new_AGEMA_signal_22072 ;
    wire new_AGEMA_signal_22073 ;
    wire new_AGEMA_signal_22074 ;
    wire new_AGEMA_signal_22075 ;
    wire new_AGEMA_signal_22076 ;
    wire new_AGEMA_signal_22077 ;
    wire new_AGEMA_signal_22078 ;
    wire new_AGEMA_signal_22079 ;
    wire new_AGEMA_signal_22080 ;
    wire new_AGEMA_signal_22081 ;
    wire new_AGEMA_signal_22082 ;
    wire new_AGEMA_signal_22083 ;
    wire new_AGEMA_signal_22084 ;
    wire new_AGEMA_signal_22085 ;
    wire new_AGEMA_signal_22086 ;
    wire new_AGEMA_signal_22087 ;
    wire new_AGEMA_signal_22088 ;
    wire new_AGEMA_signal_22089 ;
    wire new_AGEMA_signal_22090 ;
    wire new_AGEMA_signal_22091 ;
    wire new_AGEMA_signal_22092 ;
    wire new_AGEMA_signal_22093 ;
    wire new_AGEMA_signal_22094 ;
    wire new_AGEMA_signal_22095 ;
    wire new_AGEMA_signal_22096 ;
    wire new_AGEMA_signal_22097 ;
    wire new_AGEMA_signal_22098 ;
    wire new_AGEMA_signal_22099 ;
    wire new_AGEMA_signal_22100 ;
    wire new_AGEMA_signal_22101 ;
    wire new_AGEMA_signal_22102 ;
    wire new_AGEMA_signal_22103 ;
    wire new_AGEMA_signal_22104 ;
    wire new_AGEMA_signal_22105 ;
    wire new_AGEMA_signal_22106 ;
    wire new_AGEMA_signal_22107 ;
    wire new_AGEMA_signal_22108 ;
    wire new_AGEMA_signal_22109 ;
    wire new_AGEMA_signal_22110 ;
    wire new_AGEMA_signal_22111 ;
    wire new_AGEMA_signal_22112 ;
    wire new_AGEMA_signal_22113 ;
    wire new_AGEMA_signal_22114 ;
    wire new_AGEMA_signal_22115 ;
    wire new_AGEMA_signal_22116 ;
    wire new_AGEMA_signal_22117 ;
    wire new_AGEMA_signal_22118 ;
    wire new_AGEMA_signal_22119 ;
    wire new_AGEMA_signal_22120 ;
    wire new_AGEMA_signal_22121 ;
    wire new_AGEMA_signal_22122 ;
    wire new_AGEMA_signal_22123 ;
    wire new_AGEMA_signal_22124 ;
    wire new_AGEMA_signal_22125 ;
    wire new_AGEMA_signal_22126 ;
    wire new_AGEMA_signal_22127 ;
    wire new_AGEMA_signal_22128 ;
    wire new_AGEMA_signal_22129 ;
    wire new_AGEMA_signal_22130 ;
    wire new_AGEMA_signal_22131 ;
    wire new_AGEMA_signal_22132 ;
    wire new_AGEMA_signal_22133 ;
    wire new_AGEMA_signal_22134 ;
    wire new_AGEMA_signal_22135 ;
    wire new_AGEMA_signal_22136 ;
    wire new_AGEMA_signal_22137 ;
    wire new_AGEMA_signal_22138 ;
    wire new_AGEMA_signal_22139 ;
    wire new_AGEMA_signal_22140 ;
    wire new_AGEMA_signal_22141 ;
    wire new_AGEMA_signal_22142 ;
    wire new_AGEMA_signal_22143 ;
    wire new_AGEMA_signal_22144 ;
    wire new_AGEMA_signal_22145 ;
    wire new_AGEMA_signal_22146 ;
    wire new_AGEMA_signal_22147 ;
    wire new_AGEMA_signal_22148 ;
    wire new_AGEMA_signal_22149 ;
    wire new_AGEMA_signal_22150 ;
    wire new_AGEMA_signal_22151 ;
    wire new_AGEMA_signal_22152 ;
    wire new_AGEMA_signal_22153 ;
    wire new_AGEMA_signal_22154 ;
    wire new_AGEMA_signal_22155 ;
    wire new_AGEMA_signal_22156 ;
    wire new_AGEMA_signal_22157 ;
    wire new_AGEMA_signal_22158 ;
    wire new_AGEMA_signal_22159 ;
    wire new_AGEMA_signal_22160 ;
    wire new_AGEMA_signal_22161 ;
    wire new_AGEMA_signal_22162 ;
    wire new_AGEMA_signal_22163 ;
    wire new_AGEMA_signal_22164 ;
    wire new_AGEMA_signal_22165 ;
    wire new_AGEMA_signal_22166 ;
    wire new_AGEMA_signal_22167 ;
    wire new_AGEMA_signal_22168 ;
    wire new_AGEMA_signal_22169 ;
    wire new_AGEMA_signal_22170 ;
    wire new_AGEMA_signal_22171 ;
    wire new_AGEMA_signal_22172 ;
    wire new_AGEMA_signal_22173 ;
    wire new_AGEMA_signal_22174 ;
    wire new_AGEMA_signal_22175 ;
    wire new_AGEMA_signal_22176 ;
    wire new_AGEMA_signal_22177 ;
    wire new_AGEMA_signal_22178 ;
    wire new_AGEMA_signal_22179 ;
    wire new_AGEMA_signal_22180 ;
    wire new_AGEMA_signal_22181 ;
    wire new_AGEMA_signal_22182 ;
    wire new_AGEMA_signal_22183 ;
    wire new_AGEMA_signal_22184 ;
    wire new_AGEMA_signal_22185 ;
    wire new_AGEMA_signal_22186 ;
    wire new_AGEMA_signal_22187 ;
    wire new_AGEMA_signal_22188 ;
    wire new_AGEMA_signal_22189 ;
    wire new_AGEMA_signal_22190 ;
    wire new_AGEMA_signal_22191 ;
    wire new_AGEMA_signal_22192 ;
    wire new_AGEMA_signal_22193 ;
    wire new_AGEMA_signal_22194 ;
    wire new_AGEMA_signal_22195 ;
    wire new_AGEMA_signal_22196 ;
    wire new_AGEMA_signal_22197 ;
    wire new_AGEMA_signal_22198 ;
    wire new_AGEMA_signal_22199 ;
    wire new_AGEMA_signal_22200 ;
    wire new_AGEMA_signal_22201 ;
    wire new_AGEMA_signal_22202 ;
    wire new_AGEMA_signal_22203 ;
    wire new_AGEMA_signal_22204 ;
    wire new_AGEMA_signal_22205 ;
    wire new_AGEMA_signal_22206 ;
    wire new_AGEMA_signal_22207 ;
    wire new_AGEMA_signal_22208 ;
    wire new_AGEMA_signal_22209 ;
    wire new_AGEMA_signal_22210 ;
    wire new_AGEMA_signal_22211 ;
    wire new_AGEMA_signal_22212 ;
    wire new_AGEMA_signal_22213 ;
    wire new_AGEMA_signal_22214 ;
    wire new_AGEMA_signal_22215 ;
    wire new_AGEMA_signal_22216 ;
    wire new_AGEMA_signal_22217 ;
    wire new_AGEMA_signal_22218 ;
    wire new_AGEMA_signal_22219 ;
    wire new_AGEMA_signal_22220 ;
    wire new_AGEMA_signal_22221 ;
    wire new_AGEMA_signal_22222 ;
    wire new_AGEMA_signal_22223 ;
    wire new_AGEMA_signal_22224 ;
    wire new_AGEMA_signal_22225 ;
    wire new_AGEMA_signal_22226 ;
    wire new_AGEMA_signal_22227 ;
    wire new_AGEMA_signal_22228 ;
    wire new_AGEMA_signal_22229 ;
    wire new_AGEMA_signal_22230 ;
    wire new_AGEMA_signal_22231 ;
    wire new_AGEMA_signal_22232 ;
    wire new_AGEMA_signal_22233 ;
    wire new_AGEMA_signal_22234 ;
    wire new_AGEMA_signal_22235 ;
    wire new_AGEMA_signal_22236 ;
    wire new_AGEMA_signal_22237 ;
    wire new_AGEMA_signal_22238 ;
    wire new_AGEMA_signal_22239 ;
    wire new_AGEMA_signal_22240 ;
    wire new_AGEMA_signal_22241 ;
    wire new_AGEMA_signal_22242 ;
    wire new_AGEMA_signal_22243 ;
    wire new_AGEMA_signal_22244 ;
    wire new_AGEMA_signal_22245 ;
    wire new_AGEMA_signal_22246 ;
    wire new_AGEMA_signal_22247 ;
    wire new_AGEMA_signal_22248 ;
    wire new_AGEMA_signal_22249 ;
    wire new_AGEMA_signal_22250 ;
    wire new_AGEMA_signal_22251 ;
    wire new_AGEMA_signal_22252 ;
    wire new_AGEMA_signal_22253 ;
    wire new_AGEMA_signal_22254 ;
    wire new_AGEMA_signal_22255 ;
    wire new_AGEMA_signal_22256 ;
    wire new_AGEMA_signal_22257 ;
    wire new_AGEMA_signal_22258 ;
    wire new_AGEMA_signal_22259 ;
    wire new_AGEMA_signal_22260 ;
    wire new_AGEMA_signal_22261 ;
    wire new_AGEMA_signal_22262 ;
    wire new_AGEMA_signal_22263 ;
    wire new_AGEMA_signal_22264 ;
    wire new_AGEMA_signal_22265 ;
    wire new_AGEMA_signal_22266 ;
    wire new_AGEMA_signal_22267 ;
    wire new_AGEMA_signal_22268 ;
    wire new_AGEMA_signal_22269 ;
    wire new_AGEMA_signal_22270 ;
    wire new_AGEMA_signal_22271 ;
    wire new_AGEMA_signal_22272 ;
    wire new_AGEMA_signal_22273 ;
    wire new_AGEMA_signal_22274 ;
    wire new_AGEMA_signal_22275 ;
    wire new_AGEMA_signal_22276 ;
    wire new_AGEMA_signal_22277 ;
    wire new_AGEMA_signal_22278 ;
    wire new_AGEMA_signal_22279 ;
    wire new_AGEMA_signal_22280 ;
    wire new_AGEMA_signal_22281 ;
    wire new_AGEMA_signal_22282 ;
    wire new_AGEMA_signal_22283 ;
    wire new_AGEMA_signal_22284 ;
    wire new_AGEMA_signal_22285 ;
    wire new_AGEMA_signal_22286 ;
    wire new_AGEMA_signal_22287 ;
    wire new_AGEMA_signal_22288 ;
    wire new_AGEMA_signal_22289 ;
    wire new_AGEMA_signal_22290 ;
    wire new_AGEMA_signal_22291 ;
    wire new_AGEMA_signal_22292 ;
    wire new_AGEMA_signal_22293 ;
    wire new_AGEMA_signal_22294 ;
    wire new_AGEMA_signal_22295 ;
    wire new_AGEMA_signal_22296 ;
    wire new_AGEMA_signal_22297 ;
    wire new_AGEMA_signal_22298 ;
    wire new_AGEMA_signal_22299 ;
    wire new_AGEMA_signal_22300 ;
    wire new_AGEMA_signal_22301 ;
    wire new_AGEMA_signal_22302 ;
    wire new_AGEMA_signal_22303 ;
    wire new_AGEMA_signal_22304 ;
    wire new_AGEMA_signal_22305 ;
    wire new_AGEMA_signal_22306 ;
    wire new_AGEMA_signal_22307 ;
    wire new_AGEMA_signal_22308 ;
    wire new_AGEMA_signal_22309 ;
    wire new_AGEMA_signal_22310 ;
    wire new_AGEMA_signal_22311 ;
    wire new_AGEMA_signal_22312 ;
    wire new_AGEMA_signal_22313 ;
    wire new_AGEMA_signal_22314 ;
    wire new_AGEMA_signal_22315 ;
    wire new_AGEMA_signal_22316 ;
    wire new_AGEMA_signal_22317 ;
    wire new_AGEMA_signal_22318 ;
    wire new_AGEMA_signal_22319 ;
    wire new_AGEMA_signal_22320 ;
    wire new_AGEMA_signal_22321 ;
    wire new_AGEMA_signal_22322 ;
    wire new_AGEMA_signal_22323 ;
    wire new_AGEMA_signal_22324 ;
    wire new_AGEMA_signal_22325 ;
    wire new_AGEMA_signal_22326 ;
    wire new_AGEMA_signal_22327 ;
    wire new_AGEMA_signal_22328 ;
    wire new_AGEMA_signal_22329 ;
    wire new_AGEMA_signal_22330 ;
    wire new_AGEMA_signal_22331 ;
    wire new_AGEMA_signal_22332 ;
    wire new_AGEMA_signal_22333 ;
    wire new_AGEMA_signal_22334 ;
    wire new_AGEMA_signal_22335 ;
    wire new_AGEMA_signal_22336 ;
    wire new_AGEMA_signal_22337 ;
    wire new_AGEMA_signal_22338 ;
    wire new_AGEMA_signal_22339 ;
    wire new_AGEMA_signal_22340 ;
    wire new_AGEMA_signal_22341 ;
    wire new_AGEMA_signal_22342 ;
    wire new_AGEMA_signal_22343 ;
    wire new_AGEMA_signal_22344 ;
    wire new_AGEMA_signal_22345 ;
    wire new_AGEMA_signal_22346 ;
    wire new_AGEMA_signal_22347 ;
    wire new_AGEMA_signal_22348 ;
    wire new_AGEMA_signal_22349 ;
    wire new_AGEMA_signal_22350 ;
    wire new_AGEMA_signal_22351 ;
    wire new_AGEMA_signal_22352 ;
    wire new_AGEMA_signal_22353 ;
    wire new_AGEMA_signal_22354 ;
    wire new_AGEMA_signal_22355 ;
    wire new_AGEMA_signal_22356 ;
    wire new_AGEMA_signal_22357 ;
    wire new_AGEMA_signal_22358 ;
    wire new_AGEMA_signal_22359 ;
    wire new_AGEMA_signal_22360 ;
    wire new_AGEMA_signal_22361 ;
    wire new_AGEMA_signal_22362 ;
    wire new_AGEMA_signal_22363 ;
    wire new_AGEMA_signal_22364 ;
    wire new_AGEMA_signal_22365 ;
    wire new_AGEMA_signal_22366 ;
    wire new_AGEMA_signal_22367 ;
    wire new_AGEMA_signal_22368 ;
    wire new_AGEMA_signal_22369 ;
    wire new_AGEMA_signal_22370 ;
    wire new_AGEMA_signal_22371 ;
    wire new_AGEMA_signal_22372 ;
    wire new_AGEMA_signal_22373 ;
    wire new_AGEMA_signal_22374 ;
    wire new_AGEMA_signal_22375 ;
    wire new_AGEMA_signal_22376 ;
    wire new_AGEMA_signal_22377 ;
    wire new_AGEMA_signal_22378 ;
    wire new_AGEMA_signal_22379 ;
    wire new_AGEMA_signal_22380 ;
    wire new_AGEMA_signal_22381 ;
    wire new_AGEMA_signal_22382 ;
    wire new_AGEMA_signal_22383 ;
    wire new_AGEMA_signal_22384 ;
    wire new_AGEMA_signal_22385 ;
    wire new_AGEMA_signal_22386 ;
    wire new_AGEMA_signal_22387 ;
    wire new_AGEMA_signal_22388 ;
    wire new_AGEMA_signal_22389 ;
    wire new_AGEMA_signal_22390 ;
    wire new_AGEMA_signal_22391 ;
    wire new_AGEMA_signal_22392 ;
    wire new_AGEMA_signal_22393 ;
    wire new_AGEMA_signal_22394 ;
    wire new_AGEMA_signal_22395 ;
    wire new_AGEMA_signal_22396 ;
    wire new_AGEMA_signal_22397 ;
    wire new_AGEMA_signal_22398 ;
    wire new_AGEMA_signal_22399 ;
    wire new_AGEMA_signal_22400 ;
    wire new_AGEMA_signal_22401 ;
    wire new_AGEMA_signal_22402 ;
    wire new_AGEMA_signal_22403 ;
    wire new_AGEMA_signal_22404 ;
    wire new_AGEMA_signal_22405 ;
    wire new_AGEMA_signal_22406 ;
    wire new_AGEMA_signal_22407 ;
    wire new_AGEMA_signal_22408 ;
    wire new_AGEMA_signal_22409 ;
    wire new_AGEMA_signal_22410 ;
    wire new_AGEMA_signal_22411 ;
    wire new_AGEMA_signal_22412 ;
    wire new_AGEMA_signal_22413 ;
    wire new_AGEMA_signal_22414 ;
    wire new_AGEMA_signal_22415 ;
    wire new_AGEMA_signal_22416 ;
    wire new_AGEMA_signal_22417 ;
    wire new_AGEMA_signal_22418 ;
    wire new_AGEMA_signal_22419 ;
    wire new_AGEMA_signal_22420 ;
    wire new_AGEMA_signal_22421 ;
    wire new_AGEMA_signal_22422 ;
    wire new_AGEMA_signal_22423 ;
    wire new_AGEMA_signal_22424 ;
    wire new_AGEMA_signal_22425 ;
    wire new_AGEMA_signal_22426 ;
    wire new_AGEMA_signal_22427 ;
    wire new_AGEMA_signal_22428 ;
    wire new_AGEMA_signal_22429 ;
    wire new_AGEMA_signal_22430 ;
    wire new_AGEMA_signal_22431 ;
    wire new_AGEMA_signal_22432 ;
    wire new_AGEMA_signal_22433 ;
    wire new_AGEMA_signal_22434 ;
    wire new_AGEMA_signal_22435 ;
    wire new_AGEMA_signal_22436 ;
    wire new_AGEMA_signal_22437 ;
    wire new_AGEMA_signal_22438 ;
    wire new_AGEMA_signal_22439 ;
    wire new_AGEMA_signal_22440 ;
    wire new_AGEMA_signal_22441 ;
    wire new_AGEMA_signal_22442 ;
    wire new_AGEMA_signal_22443 ;
    wire new_AGEMA_signal_22444 ;
    wire new_AGEMA_signal_22445 ;
    wire new_AGEMA_signal_22446 ;
    wire new_AGEMA_signal_22447 ;
    wire new_AGEMA_signal_22448 ;
    wire new_AGEMA_signal_22449 ;
    wire new_AGEMA_signal_22450 ;
    wire new_AGEMA_signal_22451 ;
    wire new_AGEMA_signal_22452 ;
    wire new_AGEMA_signal_22453 ;
    wire new_AGEMA_signal_22454 ;
    wire new_AGEMA_signal_22455 ;
    wire new_AGEMA_signal_22456 ;
    wire new_AGEMA_signal_22457 ;
    wire new_AGEMA_signal_22458 ;
    wire new_AGEMA_signal_22459 ;
    wire new_AGEMA_signal_22460 ;
    wire new_AGEMA_signal_22461 ;
    wire new_AGEMA_signal_22462 ;
    wire new_AGEMA_signal_22463 ;
    wire new_AGEMA_signal_22464 ;
    wire new_AGEMA_signal_22465 ;
    wire new_AGEMA_signal_22466 ;
    wire new_AGEMA_signal_22467 ;
    wire new_AGEMA_signal_22468 ;
    wire new_AGEMA_signal_22469 ;
    wire new_AGEMA_signal_22470 ;
    wire new_AGEMA_signal_22471 ;
    wire new_AGEMA_signal_22472 ;
    wire new_AGEMA_signal_22473 ;
    wire new_AGEMA_signal_22474 ;
    wire new_AGEMA_signal_22475 ;
    wire new_AGEMA_signal_22476 ;
    wire new_AGEMA_signal_22477 ;
    wire new_AGEMA_signal_22478 ;
    wire new_AGEMA_signal_22479 ;
    wire new_AGEMA_signal_22480 ;
    wire new_AGEMA_signal_22481 ;
    wire new_AGEMA_signal_22482 ;
    wire new_AGEMA_signal_22483 ;
    wire new_AGEMA_signal_22484 ;
    wire new_AGEMA_signal_22485 ;
    wire new_AGEMA_signal_22486 ;
    wire new_AGEMA_signal_22487 ;
    wire new_AGEMA_signal_22488 ;
    wire new_AGEMA_signal_22489 ;
    wire new_AGEMA_signal_22490 ;
    wire new_AGEMA_signal_22491 ;
    wire new_AGEMA_signal_22492 ;
    wire new_AGEMA_signal_22493 ;
    wire new_AGEMA_signal_22494 ;
    wire new_AGEMA_signal_22495 ;
    wire new_AGEMA_signal_22496 ;
    wire new_AGEMA_signal_22497 ;
    wire new_AGEMA_signal_22498 ;
    wire new_AGEMA_signal_22499 ;
    wire new_AGEMA_signal_22500 ;
    wire new_AGEMA_signal_22501 ;
    wire new_AGEMA_signal_22502 ;
    wire new_AGEMA_signal_22503 ;
    wire new_AGEMA_signal_22504 ;
    wire new_AGEMA_signal_22505 ;
    wire new_AGEMA_signal_22506 ;
    wire new_AGEMA_signal_22507 ;
    wire new_AGEMA_signal_22508 ;
    wire new_AGEMA_signal_22509 ;
    wire new_AGEMA_signal_22510 ;
    wire new_AGEMA_signal_22511 ;
    wire new_AGEMA_signal_22512 ;
    wire new_AGEMA_signal_22513 ;
    wire new_AGEMA_signal_22514 ;
    wire new_AGEMA_signal_22515 ;
    wire new_AGEMA_signal_22516 ;
    wire new_AGEMA_signal_22517 ;
    wire new_AGEMA_signal_22518 ;
    wire new_AGEMA_signal_22519 ;
    wire new_AGEMA_signal_22520 ;
    wire new_AGEMA_signal_22521 ;
    wire new_AGEMA_signal_22522 ;
    wire new_AGEMA_signal_22523 ;
    wire new_AGEMA_signal_22524 ;
    wire new_AGEMA_signal_22525 ;
    wire new_AGEMA_signal_22526 ;
    wire new_AGEMA_signal_22527 ;
    wire new_AGEMA_signal_22528 ;
    wire new_AGEMA_signal_22529 ;
    wire new_AGEMA_signal_22530 ;
    wire new_AGEMA_signal_22531 ;
    wire new_AGEMA_signal_22532 ;
    wire new_AGEMA_signal_22533 ;
    wire new_AGEMA_signal_22534 ;
    wire new_AGEMA_signal_22535 ;
    wire new_AGEMA_signal_22536 ;
    wire new_AGEMA_signal_22537 ;
    wire new_AGEMA_signal_22538 ;
    wire new_AGEMA_signal_22539 ;
    wire new_AGEMA_signal_22540 ;
    wire new_AGEMA_signal_22541 ;
    wire new_AGEMA_signal_22542 ;
    wire new_AGEMA_signal_22543 ;
    wire new_AGEMA_signal_22544 ;
    wire new_AGEMA_signal_22545 ;
    wire new_AGEMA_signal_22546 ;
    wire new_AGEMA_signal_22547 ;
    wire new_AGEMA_signal_22548 ;
    wire new_AGEMA_signal_22549 ;
    wire new_AGEMA_signal_22550 ;
    wire new_AGEMA_signal_22551 ;
    wire new_AGEMA_signal_22552 ;
    wire new_AGEMA_signal_22553 ;
    wire new_AGEMA_signal_22554 ;
    wire new_AGEMA_signal_22555 ;
    wire new_AGEMA_signal_22556 ;
    wire new_AGEMA_signal_22557 ;
    wire new_AGEMA_signal_22558 ;
    wire new_AGEMA_signal_22559 ;
    wire new_AGEMA_signal_22560 ;
    wire new_AGEMA_signal_22561 ;
    wire new_AGEMA_signal_22562 ;
    wire new_AGEMA_signal_22563 ;
    wire new_AGEMA_signal_22564 ;
    wire new_AGEMA_signal_22565 ;
    wire new_AGEMA_signal_22566 ;
    wire new_AGEMA_signal_22567 ;
    wire new_AGEMA_signal_22568 ;
    wire new_AGEMA_signal_22569 ;
    wire new_AGEMA_signal_22570 ;
    wire new_AGEMA_signal_22571 ;
    wire new_AGEMA_signal_22572 ;
    wire new_AGEMA_signal_22573 ;
    wire new_AGEMA_signal_22574 ;
    wire new_AGEMA_signal_22575 ;
    wire new_AGEMA_signal_22576 ;
    wire new_AGEMA_signal_22577 ;
    wire new_AGEMA_signal_22578 ;
    wire new_AGEMA_signal_22579 ;
    wire new_AGEMA_signal_22580 ;
    wire new_AGEMA_signal_22581 ;
    wire new_AGEMA_signal_22582 ;
    wire new_AGEMA_signal_22583 ;
    wire new_AGEMA_signal_22584 ;
    wire new_AGEMA_signal_22585 ;
    wire new_AGEMA_signal_22586 ;
    wire new_AGEMA_signal_22587 ;
    wire new_AGEMA_signal_22588 ;
    wire new_AGEMA_signal_22589 ;
    wire new_AGEMA_signal_22590 ;
    wire new_AGEMA_signal_22591 ;
    wire new_AGEMA_signal_22592 ;
    wire new_AGEMA_signal_22593 ;
    wire new_AGEMA_signal_22594 ;
    wire new_AGEMA_signal_22595 ;
    wire new_AGEMA_signal_22596 ;
    wire new_AGEMA_signal_22597 ;
    wire new_AGEMA_signal_22598 ;
    wire new_AGEMA_signal_22599 ;
    wire new_AGEMA_signal_22600 ;
    wire new_AGEMA_signal_22601 ;
    wire new_AGEMA_signal_22602 ;
    wire new_AGEMA_signal_22603 ;
    wire new_AGEMA_signal_22604 ;
    wire new_AGEMA_signal_22605 ;
    wire new_AGEMA_signal_22606 ;
    wire new_AGEMA_signal_22607 ;
    wire new_AGEMA_signal_22608 ;
    wire new_AGEMA_signal_22609 ;
    wire new_AGEMA_signal_22610 ;
    wire new_AGEMA_signal_22611 ;
    wire new_AGEMA_signal_22612 ;
    wire new_AGEMA_signal_22613 ;
    wire new_AGEMA_signal_22614 ;
    wire new_AGEMA_signal_22615 ;
    wire new_AGEMA_signal_22616 ;
    wire new_AGEMA_signal_22617 ;
    wire new_AGEMA_signal_22618 ;
    wire new_AGEMA_signal_22619 ;
    wire new_AGEMA_signal_22620 ;
    wire new_AGEMA_signal_22621 ;
    wire new_AGEMA_signal_22622 ;
    wire new_AGEMA_signal_22623 ;
    wire new_AGEMA_signal_22624 ;
    wire new_AGEMA_signal_22625 ;
    wire new_AGEMA_signal_22626 ;
    wire new_AGEMA_signal_22627 ;
    wire new_AGEMA_signal_22628 ;
    wire new_AGEMA_signal_22629 ;
    wire new_AGEMA_signal_22630 ;
    wire new_AGEMA_signal_22631 ;
    wire new_AGEMA_signal_22632 ;
    wire new_AGEMA_signal_22633 ;
    wire new_AGEMA_signal_22634 ;
    wire new_AGEMA_signal_22635 ;
    wire new_AGEMA_signal_22636 ;
    wire new_AGEMA_signal_22637 ;
    wire new_AGEMA_signal_22638 ;
    wire new_AGEMA_signal_22639 ;
    wire new_AGEMA_signal_22640 ;
    wire new_AGEMA_signal_22641 ;
    wire new_AGEMA_signal_22642 ;
    wire new_AGEMA_signal_22643 ;
    wire new_AGEMA_signal_22644 ;
    wire new_AGEMA_signal_22645 ;
    wire new_AGEMA_signal_22646 ;
    wire new_AGEMA_signal_22647 ;
    wire new_AGEMA_signal_22648 ;
    wire new_AGEMA_signal_22649 ;
    wire new_AGEMA_signal_22650 ;
    wire new_AGEMA_signal_22651 ;
    wire new_AGEMA_signal_22652 ;
    wire new_AGEMA_signal_22653 ;
    wire new_AGEMA_signal_22654 ;
    wire new_AGEMA_signal_22655 ;
    wire new_AGEMA_signal_22656 ;
    wire new_AGEMA_signal_22657 ;
    wire new_AGEMA_signal_22658 ;
    wire new_AGEMA_signal_22659 ;
    wire new_AGEMA_signal_22660 ;
    wire new_AGEMA_signal_22661 ;
    wire new_AGEMA_signal_22662 ;
    wire new_AGEMA_signal_22663 ;
    wire new_AGEMA_signal_22664 ;
    wire new_AGEMA_signal_22665 ;
    wire new_AGEMA_signal_22666 ;
    wire new_AGEMA_signal_22667 ;
    wire new_AGEMA_signal_22668 ;
    wire new_AGEMA_signal_22669 ;
    wire new_AGEMA_signal_22670 ;
    wire new_AGEMA_signal_22671 ;
    wire new_AGEMA_signal_22672 ;
    wire new_AGEMA_signal_22673 ;
    wire new_AGEMA_signal_22674 ;
    wire new_AGEMA_signal_22675 ;
    wire new_AGEMA_signal_22676 ;
    wire new_AGEMA_signal_22677 ;
    wire new_AGEMA_signal_22678 ;
    wire new_AGEMA_signal_22679 ;
    wire new_AGEMA_signal_22680 ;
    wire new_AGEMA_signal_22681 ;
    wire new_AGEMA_signal_22682 ;
    wire new_AGEMA_signal_22683 ;
    wire new_AGEMA_signal_22684 ;
    wire new_AGEMA_signal_22685 ;
    wire new_AGEMA_signal_22686 ;
    wire new_AGEMA_signal_22687 ;
    wire new_AGEMA_signal_22688 ;
    wire new_AGEMA_signal_22689 ;
    wire new_AGEMA_signal_22690 ;
    wire new_AGEMA_signal_22691 ;
    wire new_AGEMA_signal_22692 ;
    wire new_AGEMA_signal_22693 ;
    wire new_AGEMA_signal_22694 ;
    wire new_AGEMA_signal_22695 ;
    wire new_AGEMA_signal_22696 ;
    wire new_AGEMA_signal_22697 ;
    wire new_AGEMA_signal_22698 ;
    wire new_AGEMA_signal_22699 ;
    wire new_AGEMA_signal_22700 ;
    wire new_AGEMA_signal_22701 ;
    wire new_AGEMA_signal_22702 ;
    wire new_AGEMA_signal_22703 ;
    wire new_AGEMA_signal_22704 ;
    wire new_AGEMA_signal_22705 ;
    wire new_AGEMA_signal_22706 ;
    wire new_AGEMA_signal_22707 ;
    wire new_AGEMA_signal_22708 ;
    wire new_AGEMA_signal_22709 ;
    wire new_AGEMA_signal_22710 ;
    wire new_AGEMA_signal_22711 ;
    wire new_AGEMA_signal_22712 ;
    wire new_AGEMA_signal_22713 ;
    wire new_AGEMA_signal_22714 ;
    wire new_AGEMA_signal_22715 ;
    wire new_AGEMA_signal_22716 ;
    wire new_AGEMA_signal_22717 ;
    wire new_AGEMA_signal_22718 ;
    wire new_AGEMA_signal_22719 ;
    wire new_AGEMA_signal_22720 ;
    wire new_AGEMA_signal_22721 ;
    wire new_AGEMA_signal_22722 ;
    wire new_AGEMA_signal_22723 ;
    wire new_AGEMA_signal_22724 ;
    wire new_AGEMA_signal_22725 ;
    wire new_AGEMA_signal_22726 ;
    wire new_AGEMA_signal_22727 ;
    wire new_AGEMA_signal_22728 ;
    wire new_AGEMA_signal_22729 ;
    wire new_AGEMA_signal_22730 ;
    wire new_AGEMA_signal_22731 ;
    wire new_AGEMA_signal_22732 ;
    wire new_AGEMA_signal_22733 ;
    wire new_AGEMA_signal_22734 ;
    wire new_AGEMA_signal_22735 ;
    wire new_AGEMA_signal_22736 ;
    wire new_AGEMA_signal_22737 ;
    wire new_AGEMA_signal_22738 ;
    wire new_AGEMA_signal_22739 ;
    wire new_AGEMA_signal_22740 ;
    wire new_AGEMA_signal_22741 ;
    wire new_AGEMA_signal_22742 ;
    wire new_AGEMA_signal_22743 ;
    wire new_AGEMA_signal_22744 ;
    wire new_AGEMA_signal_22745 ;
    wire new_AGEMA_signal_22746 ;
    wire new_AGEMA_signal_22747 ;
    wire new_AGEMA_signal_22748 ;
    wire new_AGEMA_signal_22749 ;
    wire new_AGEMA_signal_22750 ;
    wire new_AGEMA_signal_22751 ;
    wire new_AGEMA_signal_22752 ;
    wire new_AGEMA_signal_22753 ;
    wire new_AGEMA_signal_22754 ;
    wire new_AGEMA_signal_22755 ;
    wire new_AGEMA_signal_22756 ;
    wire new_AGEMA_signal_22757 ;
    wire new_AGEMA_signal_22758 ;
    wire new_AGEMA_signal_22759 ;
    wire new_AGEMA_signal_22760 ;
    wire new_AGEMA_signal_22761 ;
    wire new_AGEMA_signal_22762 ;
    wire new_AGEMA_signal_22763 ;
    wire new_AGEMA_signal_22764 ;
    wire new_AGEMA_signal_22765 ;
    wire new_AGEMA_signal_22766 ;
    wire new_AGEMA_signal_22767 ;
    wire new_AGEMA_signal_22768 ;
    wire new_AGEMA_signal_22769 ;
    wire new_AGEMA_signal_22770 ;
    wire new_AGEMA_signal_22771 ;
    wire new_AGEMA_signal_22772 ;
    wire new_AGEMA_signal_22773 ;
    wire new_AGEMA_signal_22774 ;
    wire new_AGEMA_signal_22775 ;
    wire new_AGEMA_signal_22776 ;
    wire new_AGEMA_signal_22777 ;
    wire new_AGEMA_signal_22778 ;
    wire new_AGEMA_signal_22779 ;
    wire new_AGEMA_signal_22780 ;
    wire new_AGEMA_signal_22781 ;
    wire new_AGEMA_signal_22782 ;
    wire new_AGEMA_signal_22783 ;
    wire new_AGEMA_signal_22784 ;
    wire new_AGEMA_signal_22785 ;
    wire new_AGEMA_signal_22786 ;
    wire new_AGEMA_signal_22787 ;
    wire new_AGEMA_signal_22788 ;
    wire new_AGEMA_signal_22789 ;
    wire new_AGEMA_signal_22790 ;
    wire new_AGEMA_signal_22791 ;
    wire new_AGEMA_signal_22792 ;
    wire new_AGEMA_signal_22793 ;
    wire new_AGEMA_signal_22794 ;
    wire new_AGEMA_signal_22795 ;
    wire new_AGEMA_signal_22796 ;
    wire new_AGEMA_signal_22797 ;
    wire new_AGEMA_signal_22798 ;
    wire new_AGEMA_signal_22799 ;
    wire new_AGEMA_signal_22800 ;
    wire new_AGEMA_signal_22801 ;
    wire new_AGEMA_signal_22802 ;
    wire new_AGEMA_signal_22803 ;
    wire new_AGEMA_signal_22804 ;
    wire new_AGEMA_signal_22805 ;
    wire new_AGEMA_signal_22806 ;
    wire new_AGEMA_signal_22807 ;
    wire new_AGEMA_signal_22808 ;
    wire new_AGEMA_signal_22809 ;
    wire new_AGEMA_signal_22810 ;
    wire new_AGEMA_signal_22811 ;
    wire new_AGEMA_signal_22812 ;
    wire new_AGEMA_signal_22813 ;
    wire new_AGEMA_signal_22814 ;
    wire new_AGEMA_signal_22815 ;
    wire new_AGEMA_signal_22816 ;
    wire new_AGEMA_signal_22817 ;
    wire new_AGEMA_signal_22818 ;
    wire new_AGEMA_signal_22819 ;
    wire new_AGEMA_signal_22820 ;
    wire new_AGEMA_signal_22821 ;
    wire new_AGEMA_signal_22822 ;
    wire new_AGEMA_signal_22823 ;
    wire new_AGEMA_signal_22824 ;
    wire new_AGEMA_signal_22825 ;
    wire new_AGEMA_signal_22826 ;
    wire new_AGEMA_signal_22827 ;
    wire new_AGEMA_signal_22828 ;
    wire new_AGEMA_signal_22829 ;
    wire new_AGEMA_signal_22830 ;
    wire new_AGEMA_signal_22831 ;
    wire new_AGEMA_signal_22832 ;
    wire new_AGEMA_signal_22833 ;
    wire new_AGEMA_signal_22834 ;
    wire new_AGEMA_signal_22835 ;
    wire new_AGEMA_signal_22836 ;
    wire new_AGEMA_signal_22837 ;
    wire new_AGEMA_signal_22838 ;
    wire new_AGEMA_signal_22839 ;
    wire new_AGEMA_signal_22840 ;
    wire new_AGEMA_signal_22841 ;
    wire new_AGEMA_signal_22842 ;
    wire new_AGEMA_signal_22843 ;
    wire new_AGEMA_signal_22844 ;
    wire new_AGEMA_signal_22845 ;
    wire new_AGEMA_signal_22846 ;
    wire new_AGEMA_signal_22847 ;
    wire new_AGEMA_signal_22848 ;
    wire new_AGEMA_signal_22849 ;
    wire new_AGEMA_signal_22850 ;
    wire new_AGEMA_signal_22851 ;
    wire new_AGEMA_signal_22852 ;
    wire new_AGEMA_signal_22853 ;
    wire new_AGEMA_signal_22854 ;
    wire new_AGEMA_signal_22855 ;
    wire new_AGEMA_signal_22856 ;
    wire new_AGEMA_signal_22857 ;
    wire new_AGEMA_signal_22858 ;
    wire new_AGEMA_signal_22859 ;
    wire new_AGEMA_signal_22860 ;
    wire new_AGEMA_signal_22861 ;
    wire new_AGEMA_signal_22862 ;
    wire new_AGEMA_signal_22863 ;
    wire new_AGEMA_signal_22864 ;
    wire new_AGEMA_signal_22865 ;
    wire new_AGEMA_signal_22866 ;
    wire new_AGEMA_signal_22867 ;
    wire new_AGEMA_signal_22868 ;
    wire new_AGEMA_signal_22869 ;
    wire new_AGEMA_signal_22870 ;
    wire new_AGEMA_signal_22871 ;
    wire new_AGEMA_signal_22872 ;
    wire new_AGEMA_signal_22873 ;
    wire new_AGEMA_signal_22874 ;
    wire new_AGEMA_signal_22875 ;
    wire new_AGEMA_signal_22876 ;
    wire new_AGEMA_signal_22877 ;
    wire new_AGEMA_signal_22878 ;
    wire new_AGEMA_signal_22879 ;
    wire new_AGEMA_signal_22880 ;
    wire new_AGEMA_signal_22881 ;
    wire new_AGEMA_signal_22882 ;
    wire new_AGEMA_signal_22883 ;
    wire new_AGEMA_signal_22884 ;
    wire new_AGEMA_signal_22885 ;
    wire new_AGEMA_signal_22886 ;
    wire new_AGEMA_signal_22887 ;
    wire new_AGEMA_signal_22888 ;
    wire new_AGEMA_signal_22889 ;
    wire new_AGEMA_signal_22890 ;
    wire new_AGEMA_signal_22891 ;
    wire new_AGEMA_signal_22892 ;
    wire new_AGEMA_signal_22893 ;
    wire new_AGEMA_signal_22894 ;
    wire new_AGEMA_signal_22895 ;
    wire new_AGEMA_signal_22896 ;
    wire new_AGEMA_signal_22897 ;
    wire new_AGEMA_signal_22898 ;
    wire new_AGEMA_signal_22899 ;
    wire new_AGEMA_signal_22900 ;
    wire new_AGEMA_signal_22901 ;
    wire new_AGEMA_signal_22902 ;
    wire new_AGEMA_signal_22903 ;
    wire new_AGEMA_signal_22904 ;
    wire new_AGEMA_signal_22905 ;
    wire new_AGEMA_signal_22906 ;
    wire new_AGEMA_signal_22907 ;
    wire new_AGEMA_signal_22908 ;
    wire new_AGEMA_signal_22909 ;
    wire new_AGEMA_signal_22910 ;
    wire new_AGEMA_signal_22911 ;
    wire new_AGEMA_signal_22912 ;
    wire new_AGEMA_signal_22913 ;
    wire new_AGEMA_signal_22914 ;
    wire new_AGEMA_signal_22915 ;
    wire new_AGEMA_signal_22916 ;
    wire new_AGEMA_signal_22917 ;
    wire new_AGEMA_signal_22918 ;
    wire new_AGEMA_signal_22919 ;
    wire new_AGEMA_signal_22920 ;
    wire new_AGEMA_signal_22921 ;
    wire new_AGEMA_signal_22922 ;
    wire new_AGEMA_signal_22923 ;
    wire new_AGEMA_signal_22924 ;
    wire new_AGEMA_signal_22925 ;
    wire new_AGEMA_signal_22926 ;
    wire new_AGEMA_signal_22927 ;
    wire new_AGEMA_signal_22928 ;
    wire new_AGEMA_signal_22929 ;
    wire new_AGEMA_signal_22930 ;
    wire new_AGEMA_signal_22931 ;
    wire new_AGEMA_signal_22932 ;
    wire new_AGEMA_signal_22933 ;
    wire new_AGEMA_signal_22934 ;
    wire new_AGEMA_signal_22935 ;
    wire new_AGEMA_signal_22936 ;
    wire new_AGEMA_signal_22937 ;
    wire new_AGEMA_signal_22938 ;
    wire new_AGEMA_signal_22939 ;
    wire new_AGEMA_signal_22940 ;
    wire new_AGEMA_signal_22941 ;
    wire new_AGEMA_signal_22942 ;
    wire new_AGEMA_signal_22943 ;
    wire new_AGEMA_signal_22944 ;
    wire new_AGEMA_signal_22945 ;
    wire new_AGEMA_signal_22946 ;
    wire new_AGEMA_signal_22947 ;
    wire new_AGEMA_signal_22948 ;
    wire new_AGEMA_signal_22949 ;
    wire new_AGEMA_signal_22950 ;
    wire new_AGEMA_signal_22951 ;
    wire new_AGEMA_signal_22952 ;
    wire new_AGEMA_signal_22953 ;
    wire new_AGEMA_signal_22954 ;
    wire new_AGEMA_signal_22955 ;
    wire new_AGEMA_signal_22956 ;
    wire new_AGEMA_signal_22957 ;
    wire new_AGEMA_signal_22958 ;
    wire new_AGEMA_signal_22959 ;
    wire new_AGEMA_signal_22960 ;
    wire new_AGEMA_signal_22961 ;
    wire new_AGEMA_signal_22962 ;
    wire new_AGEMA_signal_22963 ;
    wire new_AGEMA_signal_22964 ;
    wire new_AGEMA_signal_22965 ;
    wire new_AGEMA_signal_22966 ;
    wire new_AGEMA_signal_22967 ;
    wire new_AGEMA_signal_22968 ;
    wire new_AGEMA_signal_22969 ;
    wire new_AGEMA_signal_22970 ;
    wire new_AGEMA_signal_22971 ;
    wire new_AGEMA_signal_22972 ;
    wire new_AGEMA_signal_22973 ;
    wire new_AGEMA_signal_22974 ;
    wire new_AGEMA_signal_22975 ;
    wire new_AGEMA_signal_22976 ;
    wire new_AGEMA_signal_22977 ;
    wire new_AGEMA_signal_22978 ;
    wire new_AGEMA_signal_22979 ;
    wire new_AGEMA_signal_22980 ;
    wire new_AGEMA_signal_22981 ;
    wire new_AGEMA_signal_22982 ;
    wire new_AGEMA_signal_22983 ;
    wire new_AGEMA_signal_22984 ;
    wire new_AGEMA_signal_22985 ;
    wire new_AGEMA_signal_22986 ;
    wire new_AGEMA_signal_22987 ;
    wire new_AGEMA_signal_22988 ;
    wire new_AGEMA_signal_22989 ;
    wire new_AGEMA_signal_22990 ;
    wire new_AGEMA_signal_22991 ;
    wire new_AGEMA_signal_22992 ;
    wire new_AGEMA_signal_22993 ;
    wire new_AGEMA_signal_22994 ;
    wire new_AGEMA_signal_22995 ;
    wire new_AGEMA_signal_22996 ;
    wire new_AGEMA_signal_22997 ;
    wire new_AGEMA_signal_22998 ;
    wire new_AGEMA_signal_22999 ;
    wire new_AGEMA_signal_23000 ;
    wire new_AGEMA_signal_23001 ;
    wire new_AGEMA_signal_23002 ;
    wire new_AGEMA_signal_23003 ;
    wire new_AGEMA_signal_23004 ;
    wire new_AGEMA_signal_23005 ;
    wire new_AGEMA_signal_23006 ;
    wire new_AGEMA_signal_23007 ;
    wire new_AGEMA_signal_23008 ;
    wire new_AGEMA_signal_23009 ;
    wire new_AGEMA_signal_23010 ;
    wire new_AGEMA_signal_23011 ;
    wire new_AGEMA_signal_23012 ;
    wire new_AGEMA_signal_23013 ;
    wire new_AGEMA_signal_23014 ;
    wire new_AGEMA_signal_23015 ;
    wire new_AGEMA_signal_23016 ;
    wire new_AGEMA_signal_23017 ;
    wire new_AGEMA_signal_23018 ;
    wire new_AGEMA_signal_23019 ;
    wire new_AGEMA_signal_23020 ;
    wire new_AGEMA_signal_23021 ;
    wire new_AGEMA_signal_23022 ;
    wire new_AGEMA_signal_23023 ;
    wire new_AGEMA_signal_23024 ;
    wire new_AGEMA_signal_23025 ;
    wire new_AGEMA_signal_23026 ;
    wire new_AGEMA_signal_23027 ;
    wire new_AGEMA_signal_23028 ;
    wire new_AGEMA_signal_23029 ;
    wire new_AGEMA_signal_23030 ;
    wire new_AGEMA_signal_23031 ;
    wire new_AGEMA_signal_23032 ;
    wire new_AGEMA_signal_23033 ;
    wire new_AGEMA_signal_23034 ;
    wire new_AGEMA_signal_23035 ;
    wire new_AGEMA_signal_23036 ;
    wire new_AGEMA_signal_23037 ;
    wire new_AGEMA_signal_23038 ;
    wire new_AGEMA_signal_23039 ;
    wire new_AGEMA_signal_23040 ;
    wire new_AGEMA_signal_23041 ;
    wire new_AGEMA_signal_23042 ;
    wire new_AGEMA_signal_23043 ;
    wire new_AGEMA_signal_23044 ;
    wire new_AGEMA_signal_23045 ;
    wire new_AGEMA_signal_23046 ;
    wire new_AGEMA_signal_23047 ;
    wire new_AGEMA_signal_23048 ;
    wire new_AGEMA_signal_23049 ;
    wire new_AGEMA_signal_23050 ;
    wire new_AGEMA_signal_23051 ;
    wire new_AGEMA_signal_23052 ;
    wire new_AGEMA_signal_23053 ;
    wire new_AGEMA_signal_23054 ;
    wire new_AGEMA_signal_23055 ;
    wire new_AGEMA_signal_23056 ;
    wire new_AGEMA_signal_23057 ;
    wire new_AGEMA_signal_23058 ;
    wire new_AGEMA_signal_23059 ;
    wire new_AGEMA_signal_23060 ;
    wire new_AGEMA_signal_23061 ;
    wire new_AGEMA_signal_23062 ;
    wire new_AGEMA_signal_23063 ;
    wire new_AGEMA_signal_23064 ;
    wire new_AGEMA_signal_23065 ;
    wire new_AGEMA_signal_23066 ;
    wire new_AGEMA_signal_23067 ;
    wire new_AGEMA_signal_23068 ;
    wire new_AGEMA_signal_23069 ;
    wire new_AGEMA_signal_23070 ;
    wire new_AGEMA_signal_23071 ;
    wire new_AGEMA_signal_23072 ;
    wire new_AGEMA_signal_23073 ;
    wire new_AGEMA_signal_23074 ;
    wire new_AGEMA_signal_23075 ;
    wire new_AGEMA_signal_23076 ;
    wire new_AGEMA_signal_23077 ;
    wire new_AGEMA_signal_23078 ;
    wire new_AGEMA_signal_23079 ;
    wire new_AGEMA_signal_23080 ;
    wire new_AGEMA_signal_23081 ;
    wire new_AGEMA_signal_23082 ;
    wire new_AGEMA_signal_23083 ;
    wire new_AGEMA_signal_23084 ;
    wire new_AGEMA_signal_23085 ;
    wire new_AGEMA_signal_23086 ;
    wire new_AGEMA_signal_23087 ;
    wire new_AGEMA_signal_23088 ;
    wire new_AGEMA_signal_23089 ;
    wire new_AGEMA_signal_23090 ;
    wire new_AGEMA_signal_23091 ;
    wire new_AGEMA_signal_23092 ;
    wire new_AGEMA_signal_23093 ;
    wire new_AGEMA_signal_23094 ;
    wire new_AGEMA_signal_23095 ;
    wire new_AGEMA_signal_23096 ;
    wire new_AGEMA_signal_23097 ;
    wire new_AGEMA_signal_23098 ;
    wire new_AGEMA_signal_23099 ;
    wire new_AGEMA_signal_23100 ;
    wire new_AGEMA_signal_23101 ;
    wire new_AGEMA_signal_23102 ;
    wire new_AGEMA_signal_23103 ;
    wire new_AGEMA_signal_23104 ;
    wire new_AGEMA_signal_23105 ;
    wire new_AGEMA_signal_23106 ;
    wire new_AGEMA_signal_23107 ;
    wire new_AGEMA_signal_23108 ;
    wire new_AGEMA_signal_23109 ;
    wire new_AGEMA_signal_23110 ;
    wire new_AGEMA_signal_23111 ;
    wire new_AGEMA_signal_23112 ;
    wire new_AGEMA_signal_23113 ;
    wire new_AGEMA_signal_23114 ;
    wire new_AGEMA_signal_23115 ;
    wire new_AGEMA_signal_23116 ;
    wire new_AGEMA_signal_23117 ;
    wire new_AGEMA_signal_23118 ;
    wire new_AGEMA_signal_23119 ;
    wire new_AGEMA_signal_23120 ;
    wire new_AGEMA_signal_23121 ;
    wire new_AGEMA_signal_23122 ;
    wire new_AGEMA_signal_23123 ;
    wire new_AGEMA_signal_23124 ;
    wire new_AGEMA_signal_23125 ;
    wire new_AGEMA_signal_23126 ;
    wire new_AGEMA_signal_23127 ;
    wire new_AGEMA_signal_23128 ;
    wire new_AGEMA_signal_23129 ;
    wire new_AGEMA_signal_23130 ;
    wire new_AGEMA_signal_23131 ;
    wire new_AGEMA_signal_23132 ;
    wire new_AGEMA_signal_23133 ;
    wire new_AGEMA_signal_23134 ;
    wire new_AGEMA_signal_23135 ;
    wire new_AGEMA_signal_23136 ;
    wire new_AGEMA_signal_23137 ;
    wire new_AGEMA_signal_23138 ;
    wire new_AGEMA_signal_23139 ;
    wire new_AGEMA_signal_23140 ;
    wire new_AGEMA_signal_23141 ;
    wire new_AGEMA_signal_23142 ;
    wire new_AGEMA_signal_23143 ;
    wire new_AGEMA_signal_23144 ;
    wire new_AGEMA_signal_23145 ;
    wire new_AGEMA_signal_23146 ;
    wire new_AGEMA_signal_23147 ;
    wire new_AGEMA_signal_23148 ;
    wire new_AGEMA_signal_23149 ;
    wire new_AGEMA_signal_23150 ;
    wire new_AGEMA_signal_23151 ;
    wire new_AGEMA_signal_23152 ;
    wire new_AGEMA_signal_23153 ;
    wire new_AGEMA_signal_23154 ;
    wire new_AGEMA_signal_23155 ;
    wire new_AGEMA_signal_23156 ;
    wire new_AGEMA_signal_23157 ;
    wire new_AGEMA_signal_23158 ;
    wire new_AGEMA_signal_23159 ;
    wire new_AGEMA_signal_23160 ;
    wire new_AGEMA_signal_23161 ;
    wire new_AGEMA_signal_23162 ;
    wire new_AGEMA_signal_23163 ;
    wire new_AGEMA_signal_23164 ;
    wire new_AGEMA_signal_23165 ;
    wire new_AGEMA_signal_23166 ;
    wire new_AGEMA_signal_23167 ;
    wire new_AGEMA_signal_23168 ;
    wire new_AGEMA_signal_23169 ;
    wire new_AGEMA_signal_23170 ;
    wire new_AGEMA_signal_23171 ;
    wire new_AGEMA_signal_23172 ;
    wire new_AGEMA_signal_23173 ;
    wire new_AGEMA_signal_23174 ;
    wire new_AGEMA_signal_23175 ;
    wire new_AGEMA_signal_23176 ;
    wire new_AGEMA_signal_23177 ;
    wire new_AGEMA_signal_23178 ;
    wire new_AGEMA_signal_23179 ;
    wire new_AGEMA_signal_23180 ;
    wire new_AGEMA_signal_23181 ;
    wire new_AGEMA_signal_23182 ;
    wire new_AGEMA_signal_23183 ;
    wire new_AGEMA_signal_23184 ;
    wire new_AGEMA_signal_23185 ;
    wire new_AGEMA_signal_23186 ;
    wire new_AGEMA_signal_23187 ;
    wire new_AGEMA_signal_23188 ;
    wire new_AGEMA_signal_23189 ;
    wire new_AGEMA_signal_23190 ;
    wire new_AGEMA_signal_23191 ;
    wire new_AGEMA_signal_23192 ;
    wire new_AGEMA_signal_23193 ;
    wire new_AGEMA_signal_23194 ;
    wire new_AGEMA_signal_23195 ;
    wire new_AGEMA_signal_23196 ;
    wire new_AGEMA_signal_23197 ;
    wire new_AGEMA_signal_23198 ;
    wire new_AGEMA_signal_23199 ;
    wire new_AGEMA_signal_23200 ;
    wire new_AGEMA_signal_23201 ;
    wire new_AGEMA_signal_23202 ;
    wire new_AGEMA_signal_23203 ;
    wire new_AGEMA_signal_23204 ;
    wire new_AGEMA_signal_23205 ;
    wire new_AGEMA_signal_23206 ;
    wire new_AGEMA_signal_23207 ;
    wire new_AGEMA_signal_23208 ;
    wire new_AGEMA_signal_23209 ;
    wire new_AGEMA_signal_23210 ;
    wire new_AGEMA_signal_23211 ;
    wire new_AGEMA_signal_23212 ;
    wire new_AGEMA_signal_23213 ;
    wire new_AGEMA_signal_23214 ;
    wire new_AGEMA_signal_23215 ;
    wire new_AGEMA_signal_23216 ;
    wire new_AGEMA_signal_23217 ;
    wire new_AGEMA_signal_23218 ;
    wire new_AGEMA_signal_23219 ;
    wire new_AGEMA_signal_23220 ;
    wire new_AGEMA_signal_23221 ;
    wire new_AGEMA_signal_23222 ;
    wire new_AGEMA_signal_23223 ;
    wire new_AGEMA_signal_23224 ;
    wire new_AGEMA_signal_23225 ;
    wire new_AGEMA_signal_23226 ;
    wire new_AGEMA_signal_23227 ;
    wire new_AGEMA_signal_23228 ;
    wire new_AGEMA_signal_23229 ;
    wire new_AGEMA_signal_23230 ;
    wire new_AGEMA_signal_23231 ;
    wire new_AGEMA_signal_23232 ;
    wire new_AGEMA_signal_23233 ;
    wire new_AGEMA_signal_23234 ;
    wire new_AGEMA_signal_23235 ;
    wire new_AGEMA_signal_23236 ;
    wire new_AGEMA_signal_23237 ;
    wire new_AGEMA_signal_23238 ;
    wire new_AGEMA_signal_23239 ;
    wire new_AGEMA_signal_23240 ;
    wire new_AGEMA_signal_23241 ;
    wire new_AGEMA_signal_23242 ;
    wire new_AGEMA_signal_23243 ;
    wire new_AGEMA_signal_23244 ;
    wire new_AGEMA_signal_23245 ;
    wire new_AGEMA_signal_23246 ;
    wire new_AGEMA_signal_23247 ;
    wire new_AGEMA_signal_23248 ;
    wire new_AGEMA_signal_23249 ;
    wire new_AGEMA_signal_23250 ;
    wire new_AGEMA_signal_23251 ;
    wire new_AGEMA_signal_23252 ;
    wire new_AGEMA_signal_23253 ;
    wire new_AGEMA_signal_23254 ;
    wire new_AGEMA_signal_23255 ;
    wire new_AGEMA_signal_23256 ;
    wire new_AGEMA_signal_23257 ;
    wire new_AGEMA_signal_23258 ;
    wire new_AGEMA_signal_23259 ;
    wire new_AGEMA_signal_23260 ;
    wire new_AGEMA_signal_23261 ;
    wire new_AGEMA_signal_23262 ;
    wire new_AGEMA_signal_23263 ;
    wire new_AGEMA_signal_23264 ;
    wire new_AGEMA_signal_23265 ;
    wire new_AGEMA_signal_23266 ;
    wire new_AGEMA_signal_23267 ;
    wire new_AGEMA_signal_23268 ;
    wire new_AGEMA_signal_23269 ;
    wire new_AGEMA_signal_23270 ;
    wire new_AGEMA_signal_23271 ;
    wire new_AGEMA_signal_23272 ;
    wire new_AGEMA_signal_23273 ;
    wire new_AGEMA_signal_23274 ;
    wire new_AGEMA_signal_23275 ;
    wire new_AGEMA_signal_23276 ;
    wire new_AGEMA_signal_23277 ;
    wire new_AGEMA_signal_23278 ;
    wire new_AGEMA_signal_23279 ;
    wire new_AGEMA_signal_23280 ;
    wire new_AGEMA_signal_23281 ;
    wire new_AGEMA_signal_23282 ;
    wire new_AGEMA_signal_23283 ;
    wire new_AGEMA_signal_23284 ;
    wire new_AGEMA_signal_23285 ;
    wire new_AGEMA_signal_23286 ;
    wire new_AGEMA_signal_23287 ;
    wire new_AGEMA_signal_23288 ;
    wire new_AGEMA_signal_23289 ;
    wire new_AGEMA_signal_23290 ;
    wire new_AGEMA_signal_23291 ;
    wire new_AGEMA_signal_23292 ;
    wire new_AGEMA_signal_23293 ;
    wire new_AGEMA_signal_23294 ;
    wire new_AGEMA_signal_23295 ;
    wire new_AGEMA_signal_23296 ;
    wire new_AGEMA_signal_23297 ;
    wire new_AGEMA_signal_23298 ;
    wire new_AGEMA_signal_23299 ;
    wire new_AGEMA_signal_23300 ;
    wire new_AGEMA_signal_23301 ;
    wire new_AGEMA_signal_23302 ;
    wire new_AGEMA_signal_23303 ;
    wire new_AGEMA_signal_23304 ;
    wire new_AGEMA_signal_23305 ;
    wire new_AGEMA_signal_23306 ;
    wire new_AGEMA_signal_23307 ;
    wire new_AGEMA_signal_23308 ;
    wire new_AGEMA_signal_23309 ;
    wire new_AGEMA_signal_23310 ;
    wire new_AGEMA_signal_23311 ;
    wire new_AGEMA_signal_23312 ;
    wire new_AGEMA_signal_23313 ;
    wire new_AGEMA_signal_23314 ;
    wire new_AGEMA_signal_23315 ;
    wire new_AGEMA_signal_23316 ;
    wire new_AGEMA_signal_23317 ;
    wire new_AGEMA_signal_23318 ;
    wire new_AGEMA_signal_23319 ;
    wire new_AGEMA_signal_23320 ;
    wire new_AGEMA_signal_23321 ;
    wire new_AGEMA_signal_23322 ;
    wire new_AGEMA_signal_23323 ;
    wire new_AGEMA_signal_23324 ;
    wire new_AGEMA_signal_23325 ;
    wire new_AGEMA_signal_23326 ;
    wire new_AGEMA_signal_23327 ;
    wire new_AGEMA_signal_23328 ;
    wire new_AGEMA_signal_23329 ;
    wire new_AGEMA_signal_23330 ;
    wire new_AGEMA_signal_23331 ;
    wire new_AGEMA_signal_23332 ;
    wire new_AGEMA_signal_23333 ;
    wire new_AGEMA_signal_23334 ;
    wire new_AGEMA_signal_23335 ;
    wire new_AGEMA_signal_23336 ;
    wire new_AGEMA_signal_23337 ;
    wire new_AGEMA_signal_23338 ;
    wire new_AGEMA_signal_23339 ;
    wire new_AGEMA_signal_23340 ;
    wire new_AGEMA_signal_23341 ;
    wire new_AGEMA_signal_23342 ;
    wire new_AGEMA_signal_23343 ;
    wire new_AGEMA_signal_23344 ;
    wire new_AGEMA_signal_23345 ;
    wire new_AGEMA_signal_23346 ;
    wire new_AGEMA_signal_23347 ;
    wire new_AGEMA_signal_23348 ;
    wire new_AGEMA_signal_23349 ;
    wire new_AGEMA_signal_23350 ;
    wire new_AGEMA_signal_23351 ;
    wire new_AGEMA_signal_23352 ;
    wire new_AGEMA_signal_23353 ;
    wire new_AGEMA_signal_23354 ;
    wire new_AGEMA_signal_23355 ;
    wire new_AGEMA_signal_23356 ;
    wire new_AGEMA_signal_23357 ;
    wire new_AGEMA_signal_23358 ;
    wire new_AGEMA_signal_23359 ;
    wire new_AGEMA_signal_23360 ;
    wire new_AGEMA_signal_23361 ;
    wire new_AGEMA_signal_23362 ;
    wire new_AGEMA_signal_23363 ;
    wire new_AGEMA_signal_23364 ;
    wire new_AGEMA_signal_23365 ;
    wire new_AGEMA_signal_23366 ;
    wire new_AGEMA_signal_23367 ;
    wire new_AGEMA_signal_23368 ;
    wire new_AGEMA_signal_23369 ;
    wire new_AGEMA_signal_23370 ;
    wire new_AGEMA_signal_23371 ;
    wire new_AGEMA_signal_23372 ;
    wire new_AGEMA_signal_23373 ;
    wire new_AGEMA_signal_23374 ;
    wire new_AGEMA_signal_23375 ;
    wire new_AGEMA_signal_23376 ;
    wire new_AGEMA_signal_23377 ;
    wire new_AGEMA_signal_23378 ;
    wire new_AGEMA_signal_23379 ;
    wire new_AGEMA_signal_23380 ;
    wire new_AGEMA_signal_23381 ;
    wire new_AGEMA_signal_23382 ;
    wire new_AGEMA_signal_23383 ;
    wire new_AGEMA_signal_23384 ;
    wire new_AGEMA_signal_23385 ;
    wire new_AGEMA_signal_23386 ;
    wire new_AGEMA_signal_23387 ;
    wire new_AGEMA_signal_23388 ;
    wire new_AGEMA_signal_23389 ;
    wire new_AGEMA_signal_23390 ;
    wire new_AGEMA_signal_23391 ;
    wire new_AGEMA_signal_23392 ;
    wire new_AGEMA_signal_23393 ;
    wire new_AGEMA_signal_23394 ;
    wire new_AGEMA_signal_23395 ;
    wire new_AGEMA_signal_23396 ;
    wire new_AGEMA_signal_23397 ;
    wire new_AGEMA_signal_23398 ;
    wire new_AGEMA_signal_23399 ;
    wire new_AGEMA_signal_23400 ;
    wire new_AGEMA_signal_23401 ;
    wire new_AGEMA_signal_23402 ;
    wire new_AGEMA_signal_23403 ;
    wire new_AGEMA_signal_23404 ;
    wire new_AGEMA_signal_23405 ;
    wire new_AGEMA_signal_23406 ;
    wire new_AGEMA_signal_23407 ;
    wire new_AGEMA_signal_23408 ;
    wire new_AGEMA_signal_23409 ;
    wire new_AGEMA_signal_23410 ;
    wire new_AGEMA_signal_23411 ;
    wire new_AGEMA_signal_23412 ;
    wire new_AGEMA_signal_23413 ;
    wire new_AGEMA_signal_23414 ;
    wire new_AGEMA_signal_23415 ;
    wire new_AGEMA_signal_23416 ;
    wire new_AGEMA_signal_23417 ;
    wire new_AGEMA_signal_23418 ;
    wire new_AGEMA_signal_23419 ;
    wire new_AGEMA_signal_23420 ;
    wire new_AGEMA_signal_23421 ;
    wire new_AGEMA_signal_23422 ;
    wire new_AGEMA_signal_23423 ;
    wire new_AGEMA_signal_23424 ;
    wire new_AGEMA_signal_23425 ;
    wire new_AGEMA_signal_23426 ;
    wire new_AGEMA_signal_23427 ;
    wire new_AGEMA_signal_23428 ;
    wire new_AGEMA_signal_23429 ;
    wire new_AGEMA_signal_23430 ;
    wire new_AGEMA_signal_23431 ;
    wire new_AGEMA_signal_23432 ;
    wire new_AGEMA_signal_23433 ;
    wire new_AGEMA_signal_23434 ;
    wire new_AGEMA_signal_23435 ;
    wire new_AGEMA_signal_23436 ;
    wire new_AGEMA_signal_23437 ;
    wire new_AGEMA_signal_23438 ;
    wire new_AGEMA_signal_23439 ;
    wire new_AGEMA_signal_23440 ;
    wire new_AGEMA_signal_23441 ;
    wire new_AGEMA_signal_23442 ;
    wire new_AGEMA_signal_23443 ;
    wire new_AGEMA_signal_23444 ;
    wire new_AGEMA_signal_23445 ;
    wire new_AGEMA_signal_23446 ;
    wire new_AGEMA_signal_23447 ;
    wire new_AGEMA_signal_23448 ;
    wire new_AGEMA_signal_23449 ;
    wire new_AGEMA_signal_23450 ;
    wire new_AGEMA_signal_23451 ;
    wire new_AGEMA_signal_23452 ;
    wire new_AGEMA_signal_23453 ;
    wire new_AGEMA_signal_23454 ;
    wire new_AGEMA_signal_23455 ;
    wire new_AGEMA_signal_23456 ;
    wire new_AGEMA_signal_23457 ;
    wire new_AGEMA_signal_23458 ;
    wire new_AGEMA_signal_23459 ;
    wire new_AGEMA_signal_23460 ;
    wire new_AGEMA_signal_23461 ;
    wire new_AGEMA_signal_23462 ;
    wire new_AGEMA_signal_23463 ;
    wire new_AGEMA_signal_23464 ;
    wire new_AGEMA_signal_23465 ;
    wire new_AGEMA_signal_23466 ;
    wire new_AGEMA_signal_23467 ;
    wire new_AGEMA_signal_23468 ;
    wire new_AGEMA_signal_23469 ;
    wire new_AGEMA_signal_23470 ;
    wire new_AGEMA_signal_23471 ;
    wire new_AGEMA_signal_23472 ;
    wire new_AGEMA_signal_23473 ;
    wire new_AGEMA_signal_23474 ;
    wire new_AGEMA_signal_23475 ;
    wire new_AGEMA_signal_23476 ;
    wire new_AGEMA_signal_23477 ;
    wire new_AGEMA_signal_23478 ;
    wire new_AGEMA_signal_23479 ;
    wire new_AGEMA_signal_23480 ;
    wire new_AGEMA_signal_23481 ;
    wire new_AGEMA_signal_23482 ;
    wire new_AGEMA_signal_23483 ;
    wire new_AGEMA_signal_23484 ;
    wire new_AGEMA_signal_23485 ;
    wire new_AGEMA_signal_23486 ;
    wire new_AGEMA_signal_23487 ;
    wire new_AGEMA_signal_23488 ;
    wire new_AGEMA_signal_23489 ;
    wire new_AGEMA_signal_23490 ;
    wire new_AGEMA_signal_23491 ;
    wire new_AGEMA_signal_23492 ;
    wire new_AGEMA_signal_23493 ;
    wire new_AGEMA_signal_23494 ;
    wire new_AGEMA_signal_23495 ;
    wire new_AGEMA_signal_23496 ;
    wire new_AGEMA_signal_23497 ;
    wire new_AGEMA_signal_23498 ;
    wire new_AGEMA_signal_23499 ;
    wire new_AGEMA_signal_23500 ;
    wire new_AGEMA_signal_23501 ;
    wire new_AGEMA_signal_23502 ;
    wire new_AGEMA_signal_23503 ;
    wire new_AGEMA_signal_23504 ;
    wire new_AGEMA_signal_23505 ;
    wire new_AGEMA_signal_23506 ;
    wire new_AGEMA_signal_23507 ;
    wire new_AGEMA_signal_23508 ;
    wire new_AGEMA_signal_23509 ;
    wire new_AGEMA_signal_23510 ;
    wire new_AGEMA_signal_23511 ;
    wire new_AGEMA_signal_23512 ;
    wire new_AGEMA_signal_23513 ;
    wire new_AGEMA_signal_23514 ;
    wire new_AGEMA_signal_23515 ;
    wire new_AGEMA_signal_23516 ;
    wire new_AGEMA_signal_23517 ;
    wire new_AGEMA_signal_23518 ;
    wire new_AGEMA_signal_23519 ;
    wire new_AGEMA_signal_23520 ;
    wire new_AGEMA_signal_23521 ;
    wire new_AGEMA_signal_23522 ;
    wire new_AGEMA_signal_23523 ;
    wire new_AGEMA_signal_23524 ;
    wire new_AGEMA_signal_23525 ;
    wire new_AGEMA_signal_23526 ;
    wire new_AGEMA_signal_23527 ;
    wire new_AGEMA_signal_23528 ;
    wire new_AGEMA_signal_23529 ;
    wire new_AGEMA_signal_23530 ;
    wire new_AGEMA_signal_23531 ;
    wire new_AGEMA_signal_23532 ;
    wire new_AGEMA_signal_23533 ;
    wire new_AGEMA_signal_23534 ;
    wire new_AGEMA_signal_23535 ;
    wire new_AGEMA_signal_23536 ;
    wire new_AGEMA_signal_23537 ;
    wire new_AGEMA_signal_23538 ;
    wire new_AGEMA_signal_23539 ;
    wire new_AGEMA_signal_23540 ;
    wire new_AGEMA_signal_23541 ;
    wire new_AGEMA_signal_23542 ;
    wire new_AGEMA_signal_23543 ;
    wire new_AGEMA_signal_23544 ;
    wire new_AGEMA_signal_23545 ;
    wire new_AGEMA_signal_23546 ;
    wire new_AGEMA_signal_23547 ;
    wire new_AGEMA_signal_23548 ;
    wire new_AGEMA_signal_23549 ;
    wire new_AGEMA_signal_23550 ;
    wire new_AGEMA_signal_23551 ;
    wire new_AGEMA_signal_23552 ;
    wire new_AGEMA_signal_23553 ;
    wire new_AGEMA_signal_23554 ;
    wire new_AGEMA_signal_23555 ;
    wire new_AGEMA_signal_23556 ;
    wire new_AGEMA_signal_23557 ;
    wire new_AGEMA_signal_23558 ;
    wire new_AGEMA_signal_23559 ;
    wire new_AGEMA_signal_23560 ;
    wire new_AGEMA_signal_23561 ;
    wire new_AGEMA_signal_23562 ;
    wire new_AGEMA_signal_23563 ;
    wire new_AGEMA_signal_23564 ;
    wire new_AGEMA_signal_23565 ;
    wire new_AGEMA_signal_23566 ;
    wire new_AGEMA_signal_23567 ;
    wire new_AGEMA_signal_23568 ;
    wire new_AGEMA_signal_23569 ;
    wire new_AGEMA_signal_23570 ;
    wire new_AGEMA_signal_23571 ;
    wire new_AGEMA_signal_23572 ;
    wire new_AGEMA_signal_23573 ;
    wire new_AGEMA_signal_23574 ;
    wire new_AGEMA_signal_23575 ;
    wire new_AGEMA_signal_23576 ;
    wire new_AGEMA_signal_23577 ;
    wire new_AGEMA_signal_23578 ;
    wire new_AGEMA_signal_23579 ;
    wire new_AGEMA_signal_23580 ;
    wire new_AGEMA_signal_23581 ;
    wire new_AGEMA_signal_23582 ;
    wire new_AGEMA_signal_23583 ;
    wire new_AGEMA_signal_23584 ;
    wire new_AGEMA_signal_23585 ;
    wire new_AGEMA_signal_23586 ;
    wire new_AGEMA_signal_23587 ;
    wire new_AGEMA_signal_23588 ;
    wire new_AGEMA_signal_23589 ;
    wire new_AGEMA_signal_23590 ;
    wire new_AGEMA_signal_23591 ;
    wire new_AGEMA_signal_23592 ;
    wire new_AGEMA_signal_23593 ;
    wire new_AGEMA_signal_23594 ;
    wire new_AGEMA_signal_23595 ;
    wire new_AGEMA_signal_23596 ;
    wire new_AGEMA_signal_23597 ;
    wire new_AGEMA_signal_23598 ;
    wire new_AGEMA_signal_23599 ;
    wire new_AGEMA_signal_23600 ;
    wire new_AGEMA_signal_23601 ;
    wire new_AGEMA_signal_23602 ;
    wire new_AGEMA_signal_23603 ;
    wire new_AGEMA_signal_23604 ;
    wire new_AGEMA_signal_23605 ;
    wire new_AGEMA_signal_23606 ;
    wire new_AGEMA_signal_23607 ;
    wire new_AGEMA_signal_23608 ;
    wire new_AGEMA_signal_23609 ;
    wire new_AGEMA_signal_23610 ;
    wire new_AGEMA_signal_23611 ;
    wire new_AGEMA_signal_23612 ;
    wire new_AGEMA_signal_23613 ;
    wire new_AGEMA_signal_23614 ;
    wire new_AGEMA_signal_23615 ;
    wire new_AGEMA_signal_23616 ;
    wire new_AGEMA_signal_23617 ;
    wire new_AGEMA_signal_23618 ;
    wire new_AGEMA_signal_23619 ;
    wire new_AGEMA_signal_23620 ;
    wire new_AGEMA_signal_23621 ;
    wire new_AGEMA_signal_23622 ;
    wire new_AGEMA_signal_23623 ;
    wire new_AGEMA_signal_23624 ;
    wire new_AGEMA_signal_23625 ;
    wire new_AGEMA_signal_23626 ;
    wire new_AGEMA_signal_23627 ;
    wire new_AGEMA_signal_23628 ;
    wire new_AGEMA_signal_23629 ;
    wire new_AGEMA_signal_23630 ;
    wire new_AGEMA_signal_23631 ;
    wire new_AGEMA_signal_23632 ;
    wire new_AGEMA_signal_23633 ;
    wire new_AGEMA_signal_23634 ;
    wire new_AGEMA_signal_23635 ;
    wire new_AGEMA_signal_23636 ;
    wire new_AGEMA_signal_23637 ;
    wire new_AGEMA_signal_23638 ;
    wire new_AGEMA_signal_23639 ;
    wire new_AGEMA_signal_23640 ;
    wire new_AGEMA_signal_23641 ;
    wire new_AGEMA_signal_23642 ;
    wire new_AGEMA_signal_23643 ;
    wire new_AGEMA_signal_23644 ;
    wire new_AGEMA_signal_23645 ;
    wire new_AGEMA_signal_23646 ;
    wire new_AGEMA_signal_23647 ;
    wire new_AGEMA_signal_23648 ;
    wire new_AGEMA_signal_23649 ;
    wire new_AGEMA_signal_23650 ;
    wire new_AGEMA_signal_23651 ;
    wire new_AGEMA_signal_23652 ;
    wire new_AGEMA_signal_23653 ;
    wire new_AGEMA_signal_23654 ;
    wire new_AGEMA_signal_23655 ;
    wire new_AGEMA_signal_23656 ;
    wire new_AGEMA_signal_23657 ;
    wire new_AGEMA_signal_23658 ;
    wire new_AGEMA_signal_23659 ;
    wire new_AGEMA_signal_23660 ;
    wire new_AGEMA_signal_23661 ;
    wire new_AGEMA_signal_23662 ;
    wire new_AGEMA_signal_23663 ;
    wire new_AGEMA_signal_23664 ;
    wire new_AGEMA_signal_23665 ;
    wire new_AGEMA_signal_23666 ;
    wire new_AGEMA_signal_23667 ;
    wire new_AGEMA_signal_23668 ;
    wire new_AGEMA_signal_23669 ;
    wire new_AGEMA_signal_23670 ;
    wire new_AGEMA_signal_23671 ;
    wire new_AGEMA_signal_23672 ;
    wire new_AGEMA_signal_23673 ;
    wire new_AGEMA_signal_23674 ;
    wire new_AGEMA_signal_23675 ;
    wire new_AGEMA_signal_23676 ;
    wire new_AGEMA_signal_23677 ;
    wire new_AGEMA_signal_23678 ;
    wire new_AGEMA_signal_23679 ;
    wire new_AGEMA_signal_23680 ;
    wire new_AGEMA_signal_23681 ;
    wire new_AGEMA_signal_23682 ;
    wire new_AGEMA_signal_23683 ;
    wire new_AGEMA_signal_23684 ;
    wire new_AGEMA_signal_23685 ;
    wire new_AGEMA_signal_23686 ;
    wire new_AGEMA_signal_23687 ;
    wire new_AGEMA_signal_23688 ;
    wire new_AGEMA_signal_23689 ;
    wire new_AGEMA_signal_23690 ;
    wire new_AGEMA_signal_23691 ;
    wire new_AGEMA_signal_23692 ;
    wire new_AGEMA_signal_23693 ;
    wire new_AGEMA_signal_23694 ;
    wire new_AGEMA_signal_23695 ;
    wire new_AGEMA_signal_23696 ;
    wire new_AGEMA_signal_23697 ;
    wire new_AGEMA_signal_23698 ;
    wire new_AGEMA_signal_23699 ;
    wire new_AGEMA_signal_23700 ;
    wire new_AGEMA_signal_23701 ;
    wire new_AGEMA_signal_23702 ;
    wire new_AGEMA_signal_23703 ;
    wire new_AGEMA_signal_23704 ;
    wire new_AGEMA_signal_23705 ;
    wire new_AGEMA_signal_23706 ;
    wire new_AGEMA_signal_23707 ;
    wire new_AGEMA_signal_23708 ;
    wire new_AGEMA_signal_23709 ;
    wire new_AGEMA_signal_23710 ;
    wire new_AGEMA_signal_23711 ;
    wire new_AGEMA_signal_23712 ;
    wire new_AGEMA_signal_23713 ;
    wire new_AGEMA_signal_23714 ;
    wire new_AGEMA_signal_23715 ;
    wire new_AGEMA_signal_23716 ;
    wire new_AGEMA_signal_23717 ;
    wire new_AGEMA_signal_23718 ;
    wire new_AGEMA_signal_23719 ;
    wire new_AGEMA_signal_23720 ;
    wire new_AGEMA_signal_23721 ;
    wire new_AGEMA_signal_23722 ;
    wire new_AGEMA_signal_23723 ;
    wire new_AGEMA_signal_23724 ;
    wire new_AGEMA_signal_23725 ;
    wire new_AGEMA_signal_23726 ;
    wire new_AGEMA_signal_23727 ;
    wire new_AGEMA_signal_23728 ;
    wire new_AGEMA_signal_23729 ;
    wire new_AGEMA_signal_23730 ;
    wire new_AGEMA_signal_23731 ;
    wire new_AGEMA_signal_23732 ;
    wire new_AGEMA_signal_23733 ;
    wire new_AGEMA_signal_23734 ;
    wire new_AGEMA_signal_23735 ;
    wire new_AGEMA_signal_23736 ;
    wire new_AGEMA_signal_23737 ;
    wire new_AGEMA_signal_23738 ;
    wire new_AGEMA_signal_23739 ;
    wire new_AGEMA_signal_23740 ;
    wire new_AGEMA_signal_23741 ;
    wire new_AGEMA_signal_23742 ;
    wire new_AGEMA_signal_23743 ;
    wire new_AGEMA_signal_23744 ;
    wire new_AGEMA_signal_23745 ;
    wire new_AGEMA_signal_23746 ;
    wire new_AGEMA_signal_23747 ;
    wire new_AGEMA_signal_23748 ;
    wire new_AGEMA_signal_23749 ;
    wire new_AGEMA_signal_23750 ;
    wire new_AGEMA_signal_23751 ;
    wire new_AGEMA_signal_23752 ;
    wire new_AGEMA_signal_23753 ;
    wire new_AGEMA_signal_23754 ;
    wire new_AGEMA_signal_23755 ;
    wire new_AGEMA_signal_23756 ;
    wire new_AGEMA_signal_23757 ;
    wire new_AGEMA_signal_23758 ;
    wire new_AGEMA_signal_23759 ;
    wire new_AGEMA_signal_23760 ;
    wire new_AGEMA_signal_23761 ;
    wire new_AGEMA_signal_23762 ;
    wire new_AGEMA_signal_23763 ;
    wire new_AGEMA_signal_23764 ;
    wire new_AGEMA_signal_23765 ;
    wire new_AGEMA_signal_23766 ;
    wire new_AGEMA_signal_23767 ;
    wire new_AGEMA_signal_23768 ;
    wire new_AGEMA_signal_23769 ;
    wire new_AGEMA_signal_23770 ;
    wire new_AGEMA_signal_23771 ;
    wire new_AGEMA_signal_23772 ;
    wire new_AGEMA_signal_23773 ;
    wire new_AGEMA_signal_23774 ;
    wire new_AGEMA_signal_23775 ;
    wire new_AGEMA_signal_23776 ;
    wire new_AGEMA_signal_23777 ;
    wire new_AGEMA_signal_23778 ;
    wire new_AGEMA_signal_23779 ;
    wire new_AGEMA_signal_23780 ;
    wire new_AGEMA_signal_23781 ;
    wire new_AGEMA_signal_23782 ;
    wire new_AGEMA_signal_23783 ;
    wire new_AGEMA_signal_23784 ;
    wire new_AGEMA_signal_23785 ;
    wire new_AGEMA_signal_23786 ;
    wire new_AGEMA_signal_23787 ;
    wire new_AGEMA_signal_23788 ;
    wire new_AGEMA_signal_23789 ;
    wire new_AGEMA_signal_23790 ;
    wire new_AGEMA_signal_23791 ;
    wire new_AGEMA_signal_23792 ;
    wire new_AGEMA_signal_23793 ;
    wire new_AGEMA_signal_23794 ;
    wire new_AGEMA_signal_23795 ;
    wire new_AGEMA_signal_23796 ;
    wire new_AGEMA_signal_23797 ;
    wire new_AGEMA_signal_23798 ;
    wire new_AGEMA_signal_23799 ;
    wire new_AGEMA_signal_23800 ;
    wire new_AGEMA_signal_23801 ;
    wire new_AGEMA_signal_23802 ;
    wire new_AGEMA_signal_23803 ;
    wire new_AGEMA_signal_23804 ;
    wire new_AGEMA_signal_23805 ;
    wire new_AGEMA_signal_23806 ;
    wire new_AGEMA_signal_23807 ;
    wire new_AGEMA_signal_23808 ;
    wire new_AGEMA_signal_23809 ;
    wire new_AGEMA_signal_23810 ;
    wire new_AGEMA_signal_23811 ;
    wire new_AGEMA_signal_23812 ;
    wire new_AGEMA_signal_23813 ;
    wire new_AGEMA_signal_23814 ;
    wire new_AGEMA_signal_23815 ;
    wire new_AGEMA_signal_23816 ;
    wire new_AGEMA_signal_23817 ;
    wire new_AGEMA_signal_23818 ;
    wire new_AGEMA_signal_23819 ;
    wire new_AGEMA_signal_23820 ;
    wire new_AGEMA_signal_23821 ;
    wire new_AGEMA_signal_23822 ;
    wire new_AGEMA_signal_23823 ;
    wire new_AGEMA_signal_23824 ;
    wire new_AGEMA_signal_23825 ;
    wire new_AGEMA_signal_23826 ;
    wire new_AGEMA_signal_23827 ;
    wire new_AGEMA_signal_23828 ;
    wire new_AGEMA_signal_23829 ;
    wire new_AGEMA_signal_23830 ;
    wire new_AGEMA_signal_23831 ;
    wire new_AGEMA_signal_23832 ;
    wire new_AGEMA_signal_23833 ;
    wire new_AGEMA_signal_23834 ;
    wire new_AGEMA_signal_23835 ;
    wire new_AGEMA_signal_23836 ;
    wire new_AGEMA_signal_23837 ;
    wire new_AGEMA_signal_23838 ;
    wire new_AGEMA_signal_23839 ;
    wire new_AGEMA_signal_23840 ;
    wire new_AGEMA_signal_23841 ;
    wire new_AGEMA_signal_23842 ;
    wire new_AGEMA_signal_23843 ;
    wire new_AGEMA_signal_23844 ;
    wire new_AGEMA_signal_23845 ;
    wire new_AGEMA_signal_23846 ;
    wire new_AGEMA_signal_23847 ;
    wire new_AGEMA_signal_23848 ;
    wire new_AGEMA_signal_23849 ;
    wire new_AGEMA_signal_23850 ;
    wire new_AGEMA_signal_23851 ;
    wire new_AGEMA_signal_23852 ;
    wire new_AGEMA_signal_23853 ;
    wire new_AGEMA_signal_23854 ;
    wire new_AGEMA_signal_23855 ;
    wire new_AGEMA_signal_23856 ;
    wire new_AGEMA_signal_23857 ;
    wire new_AGEMA_signal_23858 ;
    wire new_AGEMA_signal_23859 ;
    wire new_AGEMA_signal_23860 ;
    wire new_AGEMA_signal_23861 ;
    wire new_AGEMA_signal_23862 ;
    wire new_AGEMA_signal_23863 ;
    wire new_AGEMA_signal_23864 ;
    wire new_AGEMA_signal_23865 ;
    wire new_AGEMA_signal_23866 ;
    wire new_AGEMA_signal_23867 ;
    wire new_AGEMA_signal_23868 ;
    wire new_AGEMA_signal_23869 ;
    wire new_AGEMA_signal_23870 ;
    wire new_AGEMA_signal_23871 ;
    wire new_AGEMA_signal_23872 ;
    wire new_AGEMA_signal_23873 ;
    wire new_AGEMA_signal_23874 ;
    wire new_AGEMA_signal_23875 ;
    wire new_AGEMA_signal_23876 ;
    wire new_AGEMA_signal_23877 ;
    wire new_AGEMA_signal_23878 ;
    wire new_AGEMA_signal_23879 ;
    wire new_AGEMA_signal_23880 ;
    wire new_AGEMA_signal_23881 ;
    wire new_AGEMA_signal_23882 ;
    wire new_AGEMA_signal_23883 ;
    wire new_AGEMA_signal_23884 ;
    wire new_AGEMA_signal_23885 ;
    wire new_AGEMA_signal_23886 ;
    wire new_AGEMA_signal_23887 ;
    wire new_AGEMA_signal_23888 ;
    wire new_AGEMA_signal_23889 ;
    wire new_AGEMA_signal_23890 ;
    wire new_AGEMA_signal_23891 ;
    wire new_AGEMA_signal_23892 ;
    wire new_AGEMA_signal_23893 ;
    wire new_AGEMA_signal_23894 ;
    wire new_AGEMA_signal_23895 ;
    wire new_AGEMA_signal_23896 ;
    wire new_AGEMA_signal_23897 ;
    wire new_AGEMA_signal_23898 ;
    wire new_AGEMA_signal_23899 ;
    wire new_AGEMA_signal_23900 ;
    wire new_AGEMA_signal_23901 ;
    wire new_AGEMA_signal_23902 ;
    wire new_AGEMA_signal_23903 ;
    wire new_AGEMA_signal_23904 ;
    wire new_AGEMA_signal_23905 ;
    wire new_AGEMA_signal_23906 ;
    wire new_AGEMA_signal_23907 ;
    wire new_AGEMA_signal_23908 ;
    wire new_AGEMA_signal_23909 ;
    wire new_AGEMA_signal_23910 ;
    wire new_AGEMA_signal_23911 ;
    wire new_AGEMA_signal_23912 ;
    wire new_AGEMA_signal_23913 ;
    wire new_AGEMA_signal_23914 ;
    wire new_AGEMA_signal_23915 ;
    wire new_AGEMA_signal_23916 ;
    wire new_AGEMA_signal_23917 ;
    wire new_AGEMA_signal_23918 ;
    wire new_AGEMA_signal_23919 ;
    wire new_AGEMA_signal_23920 ;
    wire new_AGEMA_signal_23921 ;
    wire new_AGEMA_signal_23922 ;
    wire new_AGEMA_signal_23923 ;
    wire new_AGEMA_signal_23924 ;
    wire new_AGEMA_signal_23925 ;
    wire new_AGEMA_signal_23926 ;
    wire new_AGEMA_signal_23927 ;
    wire new_AGEMA_signal_23928 ;
    wire new_AGEMA_signal_23929 ;
    wire new_AGEMA_signal_23930 ;
    wire new_AGEMA_signal_23931 ;
    wire new_AGEMA_signal_23932 ;
    wire new_AGEMA_signal_23933 ;
    wire new_AGEMA_signal_23934 ;
    wire new_AGEMA_signal_23935 ;
    wire new_AGEMA_signal_23936 ;
    wire new_AGEMA_signal_23937 ;
    wire new_AGEMA_signal_23938 ;
    wire new_AGEMA_signal_23939 ;
    wire new_AGEMA_signal_23940 ;
    wire new_AGEMA_signal_23941 ;
    wire new_AGEMA_signal_23942 ;
    wire new_AGEMA_signal_23943 ;
    wire new_AGEMA_signal_23944 ;
    wire new_AGEMA_signal_23945 ;
    wire new_AGEMA_signal_23946 ;
    wire new_AGEMA_signal_23947 ;
    wire new_AGEMA_signal_23948 ;
    wire new_AGEMA_signal_23949 ;
    wire new_AGEMA_signal_23950 ;
    wire new_AGEMA_signal_23951 ;
    wire new_AGEMA_signal_23952 ;
    wire new_AGEMA_signal_23953 ;
    wire new_AGEMA_signal_23954 ;
    wire new_AGEMA_signal_23955 ;
    wire new_AGEMA_signal_23956 ;
    wire new_AGEMA_signal_23957 ;
    wire new_AGEMA_signal_23958 ;
    wire new_AGEMA_signal_23959 ;
    wire new_AGEMA_signal_23960 ;
    wire new_AGEMA_signal_23961 ;
    wire new_AGEMA_signal_23962 ;
    wire new_AGEMA_signal_23963 ;
    wire new_AGEMA_signal_23964 ;
    wire new_AGEMA_signal_23965 ;
    wire new_AGEMA_signal_23966 ;
    wire new_AGEMA_signal_23967 ;
    wire new_AGEMA_signal_23968 ;
    wire new_AGEMA_signal_23969 ;
    wire new_AGEMA_signal_23970 ;
    wire new_AGEMA_signal_23971 ;
    wire new_AGEMA_signal_23972 ;
    wire new_AGEMA_signal_23973 ;
    wire new_AGEMA_signal_23974 ;
    wire new_AGEMA_signal_23975 ;
    wire new_AGEMA_signal_23976 ;
    wire new_AGEMA_signal_23977 ;
    wire new_AGEMA_signal_23978 ;
    wire new_AGEMA_signal_23979 ;
    wire new_AGEMA_signal_23980 ;
    wire new_AGEMA_signal_23981 ;
    wire new_AGEMA_signal_23982 ;
    wire new_AGEMA_signal_23983 ;
    wire new_AGEMA_signal_23984 ;
    wire new_AGEMA_signal_23985 ;
    wire new_AGEMA_signal_23986 ;
    wire new_AGEMA_signal_23987 ;
    wire new_AGEMA_signal_23988 ;
    wire new_AGEMA_signal_23989 ;
    wire new_AGEMA_signal_23990 ;
    wire new_AGEMA_signal_23991 ;
    wire new_AGEMA_signal_23992 ;
    wire new_AGEMA_signal_23993 ;
    wire new_AGEMA_signal_23994 ;
    wire new_AGEMA_signal_23995 ;
    wire new_AGEMA_signal_23996 ;
    wire new_AGEMA_signal_23997 ;
    wire new_AGEMA_signal_23998 ;
    wire new_AGEMA_signal_23999 ;
    wire new_AGEMA_signal_24000 ;
    wire new_AGEMA_signal_24001 ;
    wire new_AGEMA_signal_24002 ;
    wire new_AGEMA_signal_24003 ;
    wire new_AGEMA_signal_24004 ;
    wire new_AGEMA_signal_24005 ;
    wire new_AGEMA_signal_24006 ;
    wire new_AGEMA_signal_24007 ;
    wire new_AGEMA_signal_24008 ;
    wire new_AGEMA_signal_24009 ;
    wire new_AGEMA_signal_24010 ;
    wire new_AGEMA_signal_24011 ;
    wire new_AGEMA_signal_24012 ;
    wire new_AGEMA_signal_24013 ;
    wire new_AGEMA_signal_24014 ;
    wire new_AGEMA_signal_24015 ;
    wire new_AGEMA_signal_24016 ;
    wire new_AGEMA_signal_24017 ;
    wire new_AGEMA_signal_24018 ;
    wire new_AGEMA_signal_24019 ;
    wire new_AGEMA_signal_24020 ;
    wire new_AGEMA_signal_24021 ;
    wire new_AGEMA_signal_24022 ;
    wire new_AGEMA_signal_24023 ;
    wire new_AGEMA_signal_24024 ;
    wire new_AGEMA_signal_24025 ;
    wire new_AGEMA_signal_24026 ;
    wire new_AGEMA_signal_24027 ;
    wire new_AGEMA_signal_24028 ;
    wire new_AGEMA_signal_24029 ;
    wire new_AGEMA_signal_24030 ;
    wire new_AGEMA_signal_24031 ;
    wire new_AGEMA_signal_24032 ;
    wire new_AGEMA_signal_24033 ;
    wire new_AGEMA_signal_24034 ;
    wire new_AGEMA_signal_24035 ;
    wire new_AGEMA_signal_24036 ;
    wire new_AGEMA_signal_24037 ;
    wire new_AGEMA_signal_24038 ;
    wire new_AGEMA_signal_24039 ;
    wire new_AGEMA_signal_24040 ;
    wire new_AGEMA_signal_24041 ;
    wire new_AGEMA_signal_24042 ;
    wire new_AGEMA_signal_24043 ;
    wire new_AGEMA_signal_24044 ;
    wire new_AGEMA_signal_24045 ;
    wire new_AGEMA_signal_24046 ;
    wire new_AGEMA_signal_24047 ;
    wire new_AGEMA_signal_24048 ;
    wire new_AGEMA_signal_24049 ;
    wire new_AGEMA_signal_24050 ;
    wire new_AGEMA_signal_24051 ;
    wire new_AGEMA_signal_24052 ;
    wire new_AGEMA_signal_24053 ;
    wire new_AGEMA_signal_24054 ;
    wire new_AGEMA_signal_24055 ;
    wire new_AGEMA_signal_24056 ;
    wire new_AGEMA_signal_24057 ;
    wire new_AGEMA_signal_24058 ;
    wire new_AGEMA_signal_24059 ;
    wire new_AGEMA_signal_24060 ;
    wire new_AGEMA_signal_24061 ;
    wire new_AGEMA_signal_24062 ;
    wire new_AGEMA_signal_24063 ;
    wire new_AGEMA_signal_24064 ;
    wire new_AGEMA_signal_24065 ;
    wire new_AGEMA_signal_24066 ;
    wire new_AGEMA_signal_24067 ;
    wire new_AGEMA_signal_24068 ;
    wire new_AGEMA_signal_24069 ;
    wire new_AGEMA_signal_24070 ;
    wire new_AGEMA_signal_24071 ;
    wire new_AGEMA_signal_24072 ;
    wire new_AGEMA_signal_24073 ;
    wire new_AGEMA_signal_24074 ;
    wire new_AGEMA_signal_24075 ;
    wire new_AGEMA_signal_24076 ;
    wire new_AGEMA_signal_24077 ;
    wire new_AGEMA_signal_24078 ;
    wire new_AGEMA_signal_24079 ;
    wire new_AGEMA_signal_24080 ;
    wire new_AGEMA_signal_24081 ;
    wire new_AGEMA_signal_24082 ;
    wire new_AGEMA_signal_24083 ;
    wire new_AGEMA_signal_24084 ;
    wire new_AGEMA_signal_24085 ;
    wire new_AGEMA_signal_24086 ;
    wire new_AGEMA_signal_24087 ;
    wire new_AGEMA_signal_24088 ;
    wire new_AGEMA_signal_24089 ;
    wire new_AGEMA_signal_24090 ;
    wire new_AGEMA_signal_24091 ;
    wire new_AGEMA_signal_24092 ;
    wire new_AGEMA_signal_24093 ;
    wire new_AGEMA_signal_24094 ;
    wire new_AGEMA_signal_24095 ;
    wire new_AGEMA_signal_24096 ;
    wire new_AGEMA_signal_24097 ;
    wire new_AGEMA_signal_24098 ;
    wire new_AGEMA_signal_24099 ;
    wire new_AGEMA_signal_24100 ;
    wire new_AGEMA_signal_24101 ;
    wire new_AGEMA_signal_24102 ;
    wire new_AGEMA_signal_24103 ;
    wire new_AGEMA_signal_24104 ;
    wire new_AGEMA_signal_24105 ;
    wire new_AGEMA_signal_24106 ;
    wire new_AGEMA_signal_24107 ;
    wire new_AGEMA_signal_24108 ;
    wire new_AGEMA_signal_24109 ;
    wire new_AGEMA_signal_24110 ;
    wire new_AGEMA_signal_24111 ;
    wire new_AGEMA_signal_24112 ;
    wire new_AGEMA_signal_24113 ;
    wire new_AGEMA_signal_24114 ;
    wire new_AGEMA_signal_24115 ;
    wire new_AGEMA_signal_24116 ;
    wire new_AGEMA_signal_24117 ;
    wire new_AGEMA_signal_24118 ;
    wire new_AGEMA_signal_24119 ;
    wire new_AGEMA_signal_24120 ;
    wire new_AGEMA_signal_24121 ;
    wire new_AGEMA_signal_24122 ;
    wire new_AGEMA_signal_24123 ;
    wire new_AGEMA_signal_24124 ;
    wire new_AGEMA_signal_24125 ;
    wire new_AGEMA_signal_24126 ;
    wire new_AGEMA_signal_24127 ;
    wire new_AGEMA_signal_24128 ;
    wire new_AGEMA_signal_24129 ;
    wire new_AGEMA_signal_24130 ;
    wire new_AGEMA_signal_24131 ;
    wire new_AGEMA_signal_24132 ;
    wire new_AGEMA_signal_24133 ;
    wire new_AGEMA_signal_24134 ;
    wire new_AGEMA_signal_24135 ;
    wire new_AGEMA_signal_24136 ;
    wire new_AGEMA_signal_24137 ;
    wire new_AGEMA_signal_24138 ;
    wire new_AGEMA_signal_24139 ;
    wire new_AGEMA_signal_24140 ;
    wire new_AGEMA_signal_24141 ;
    wire new_AGEMA_signal_24142 ;
    wire new_AGEMA_signal_24143 ;
    wire new_AGEMA_signal_24144 ;
    wire new_AGEMA_signal_24145 ;
    wire new_AGEMA_signal_24146 ;
    wire new_AGEMA_signal_24147 ;
    wire new_AGEMA_signal_24148 ;
    wire new_AGEMA_signal_24149 ;
    wire new_AGEMA_signal_24150 ;
    wire new_AGEMA_signal_24151 ;
    wire new_AGEMA_signal_24152 ;
    wire new_AGEMA_signal_24153 ;
    wire new_AGEMA_signal_24154 ;
    wire new_AGEMA_signal_24155 ;
    wire new_AGEMA_signal_24156 ;
    wire new_AGEMA_signal_24157 ;
    wire new_AGEMA_signal_24158 ;
    wire new_AGEMA_signal_24159 ;
    wire new_AGEMA_signal_24160 ;
    wire new_AGEMA_signal_24161 ;
    wire new_AGEMA_signal_24162 ;
    wire new_AGEMA_signal_24163 ;
    wire new_AGEMA_signal_24164 ;
    wire new_AGEMA_signal_24165 ;
    wire new_AGEMA_signal_24166 ;
    wire new_AGEMA_signal_24167 ;
    wire new_AGEMA_signal_24168 ;
    wire new_AGEMA_signal_24169 ;
    wire new_AGEMA_signal_24170 ;
    wire new_AGEMA_signal_24171 ;
    wire new_AGEMA_signal_24172 ;
    wire new_AGEMA_signal_24173 ;
    wire new_AGEMA_signal_24174 ;
    wire new_AGEMA_signal_24175 ;
    wire new_AGEMA_signal_24176 ;
    wire new_AGEMA_signal_24177 ;
    wire new_AGEMA_signal_24178 ;
    wire new_AGEMA_signal_24179 ;
    wire new_AGEMA_signal_24180 ;
    wire new_AGEMA_signal_24181 ;
    wire new_AGEMA_signal_24182 ;
    wire new_AGEMA_signal_24183 ;
    wire new_AGEMA_signal_24184 ;
    wire new_AGEMA_signal_24185 ;
    wire new_AGEMA_signal_24186 ;
    wire new_AGEMA_signal_24187 ;
    wire new_AGEMA_signal_24188 ;
    wire new_AGEMA_signal_24189 ;
    wire new_AGEMA_signal_24190 ;
    wire new_AGEMA_signal_24191 ;
    wire new_AGEMA_signal_24192 ;
    wire new_AGEMA_signal_24193 ;
    wire new_AGEMA_signal_24194 ;
    wire new_AGEMA_signal_24195 ;
    wire new_AGEMA_signal_24196 ;
    wire new_AGEMA_signal_24197 ;
    wire new_AGEMA_signal_24198 ;
    wire new_AGEMA_signal_24199 ;
    wire new_AGEMA_signal_24200 ;
    wire new_AGEMA_signal_24201 ;
    wire new_AGEMA_signal_24202 ;
    wire new_AGEMA_signal_24203 ;
    wire new_AGEMA_signal_24204 ;
    wire new_AGEMA_signal_24205 ;
    wire new_AGEMA_signal_24206 ;
    wire new_AGEMA_signal_24207 ;
    wire new_AGEMA_signal_24208 ;
    wire new_AGEMA_signal_24209 ;
    wire new_AGEMA_signal_24210 ;
    wire new_AGEMA_signal_24211 ;
    wire new_AGEMA_signal_24212 ;
    wire new_AGEMA_signal_24213 ;
    wire new_AGEMA_signal_24214 ;
    wire new_AGEMA_signal_24215 ;
    wire new_AGEMA_signal_24216 ;
    wire new_AGEMA_signal_24217 ;
    wire new_AGEMA_signal_24218 ;
    wire new_AGEMA_signal_24219 ;
    wire new_AGEMA_signal_24220 ;
    wire new_AGEMA_signal_24221 ;
    wire new_AGEMA_signal_24222 ;
    wire new_AGEMA_signal_24223 ;
    wire new_AGEMA_signal_24224 ;
    wire new_AGEMA_signal_24225 ;
    wire new_AGEMA_signal_24226 ;
    wire new_AGEMA_signal_24227 ;
    wire new_AGEMA_signal_24228 ;
    wire new_AGEMA_signal_24229 ;
    wire new_AGEMA_signal_24230 ;
    wire new_AGEMA_signal_24231 ;
    wire new_AGEMA_signal_24232 ;
    wire new_AGEMA_signal_24233 ;
    wire new_AGEMA_signal_24234 ;
    wire new_AGEMA_signal_24235 ;
    wire new_AGEMA_signal_24236 ;
    wire new_AGEMA_signal_24237 ;
    wire new_AGEMA_signal_24238 ;
    wire new_AGEMA_signal_24239 ;
    wire new_AGEMA_signal_24240 ;
    wire new_AGEMA_signal_24241 ;
    wire new_AGEMA_signal_24242 ;
    wire new_AGEMA_signal_24243 ;
    wire new_AGEMA_signal_24244 ;
    wire new_AGEMA_signal_24245 ;
    wire new_AGEMA_signal_24246 ;
    wire new_AGEMA_signal_24247 ;
    wire new_AGEMA_signal_24248 ;
    wire new_AGEMA_signal_24249 ;
    wire new_AGEMA_signal_24250 ;
    wire new_AGEMA_signal_24251 ;
    wire new_AGEMA_signal_24252 ;
    wire new_AGEMA_signal_24253 ;
    wire new_AGEMA_signal_24254 ;
    wire new_AGEMA_signal_24255 ;
    wire new_AGEMA_signal_24256 ;
    wire new_AGEMA_signal_24257 ;
    wire new_AGEMA_signal_24258 ;
    wire new_AGEMA_signal_24259 ;
    wire new_AGEMA_signal_24260 ;
    wire new_AGEMA_signal_24261 ;
    wire new_AGEMA_signal_24262 ;
    wire new_AGEMA_signal_24263 ;
    wire new_AGEMA_signal_24264 ;
    wire new_AGEMA_signal_24265 ;
    wire new_AGEMA_signal_24266 ;
    wire new_AGEMA_signal_24267 ;
    wire new_AGEMA_signal_24268 ;
    wire new_AGEMA_signal_24269 ;
    wire new_AGEMA_signal_24270 ;
    wire new_AGEMA_signal_24271 ;
    wire new_AGEMA_signal_24272 ;
    wire new_AGEMA_signal_24273 ;
    wire new_AGEMA_signal_24274 ;
    wire new_AGEMA_signal_24275 ;
    wire new_AGEMA_signal_24276 ;
    wire new_AGEMA_signal_24277 ;
    wire new_AGEMA_signal_24278 ;
    wire new_AGEMA_signal_24279 ;
    wire new_AGEMA_signal_24280 ;
    wire new_AGEMA_signal_24281 ;
    wire new_AGEMA_signal_24282 ;
    wire new_AGEMA_signal_24283 ;
    wire new_AGEMA_signal_24284 ;
    wire new_AGEMA_signal_24285 ;
    wire new_AGEMA_signal_24286 ;
    wire new_AGEMA_signal_24287 ;
    wire new_AGEMA_signal_24288 ;
    wire new_AGEMA_signal_24289 ;
    wire new_AGEMA_signal_24290 ;
    wire new_AGEMA_signal_24291 ;
    wire new_AGEMA_signal_24292 ;
    wire new_AGEMA_signal_24293 ;
    wire new_AGEMA_signal_24294 ;
    wire new_AGEMA_signal_24295 ;
    wire new_AGEMA_signal_24296 ;
    wire new_AGEMA_signal_24297 ;
    wire new_AGEMA_signal_24298 ;
    wire new_AGEMA_signal_24299 ;
    wire new_AGEMA_signal_24300 ;
    wire new_AGEMA_signal_24301 ;
    wire new_AGEMA_signal_24302 ;
    wire new_AGEMA_signal_24303 ;
    wire new_AGEMA_signal_24304 ;
    wire new_AGEMA_signal_24305 ;
    wire new_AGEMA_signal_24306 ;
    wire new_AGEMA_signal_24307 ;
    wire new_AGEMA_signal_24308 ;
    wire new_AGEMA_signal_24309 ;
    wire new_AGEMA_signal_24310 ;
    wire new_AGEMA_signal_24311 ;
    wire new_AGEMA_signal_24312 ;
    wire new_AGEMA_signal_24313 ;
    wire new_AGEMA_signal_24314 ;
    wire new_AGEMA_signal_24315 ;
    wire new_AGEMA_signal_24316 ;
    wire new_AGEMA_signal_24317 ;
    wire new_AGEMA_signal_24318 ;
    wire new_AGEMA_signal_24319 ;
    wire new_AGEMA_signal_24320 ;
    wire new_AGEMA_signal_24321 ;
    wire new_AGEMA_signal_24322 ;
    wire new_AGEMA_signal_24323 ;
    wire new_AGEMA_signal_24324 ;
    wire new_AGEMA_signal_24325 ;
    wire new_AGEMA_signal_24326 ;
    wire new_AGEMA_signal_24327 ;
    wire new_AGEMA_signal_24328 ;
    wire new_AGEMA_signal_24329 ;
    wire new_AGEMA_signal_24330 ;
    wire new_AGEMA_signal_24331 ;
    wire new_AGEMA_signal_24332 ;
    wire new_AGEMA_signal_24333 ;
    wire new_AGEMA_signal_24334 ;
    wire new_AGEMA_signal_24335 ;
    wire new_AGEMA_signal_24336 ;
    wire new_AGEMA_signal_24337 ;
    wire new_AGEMA_signal_24338 ;
    wire new_AGEMA_signal_24339 ;
    wire new_AGEMA_signal_24340 ;
    wire new_AGEMA_signal_24341 ;
    wire new_AGEMA_signal_24342 ;
    wire new_AGEMA_signal_24343 ;
    wire new_AGEMA_signal_24344 ;
    wire new_AGEMA_signal_24345 ;
    wire new_AGEMA_signal_24346 ;
    wire new_AGEMA_signal_24347 ;
    wire new_AGEMA_signal_24348 ;
    wire new_AGEMA_signal_24349 ;
    wire new_AGEMA_signal_24350 ;
    wire new_AGEMA_signal_24351 ;
    wire new_AGEMA_signal_24352 ;
    wire new_AGEMA_signal_24353 ;
    wire new_AGEMA_signal_24354 ;
    wire new_AGEMA_signal_24355 ;
    wire new_AGEMA_signal_24356 ;
    wire new_AGEMA_signal_24357 ;
    wire new_AGEMA_signal_24358 ;
    wire new_AGEMA_signal_24359 ;
    wire new_AGEMA_signal_24360 ;
    wire new_AGEMA_signal_24361 ;
    wire new_AGEMA_signal_24362 ;
    wire new_AGEMA_signal_24363 ;
    wire new_AGEMA_signal_24364 ;
    wire new_AGEMA_signal_24365 ;
    wire new_AGEMA_signal_24366 ;
    wire new_AGEMA_signal_24367 ;
    wire new_AGEMA_signal_24368 ;
    wire new_AGEMA_signal_24369 ;
    wire new_AGEMA_signal_24370 ;
    wire new_AGEMA_signal_24371 ;
    wire new_AGEMA_signal_24372 ;
    wire new_AGEMA_signal_24373 ;
    wire new_AGEMA_signal_24374 ;
    wire new_AGEMA_signal_24375 ;
    wire new_AGEMA_signal_24376 ;
    wire new_AGEMA_signal_24377 ;
    wire new_AGEMA_signal_24378 ;
    wire new_AGEMA_signal_24379 ;
    wire new_AGEMA_signal_24380 ;
    wire new_AGEMA_signal_24381 ;
    wire new_AGEMA_signal_24382 ;
    wire new_AGEMA_signal_24383 ;
    wire new_AGEMA_signal_24384 ;
    wire new_AGEMA_signal_24385 ;
    wire new_AGEMA_signal_24386 ;
    wire new_AGEMA_signal_24387 ;
    wire new_AGEMA_signal_24388 ;
    wire new_AGEMA_signal_24389 ;
    wire new_AGEMA_signal_24390 ;
    wire new_AGEMA_signal_24391 ;
    wire new_AGEMA_signal_24392 ;
    wire new_AGEMA_signal_24393 ;
    wire new_AGEMA_signal_24394 ;
    wire new_AGEMA_signal_24395 ;
    wire new_AGEMA_signal_24396 ;
    wire new_AGEMA_signal_24397 ;
    wire new_AGEMA_signal_24398 ;
    wire new_AGEMA_signal_24399 ;
    wire new_AGEMA_signal_24400 ;
    wire new_AGEMA_signal_24401 ;
    wire new_AGEMA_signal_24402 ;
    wire new_AGEMA_signal_24403 ;
    wire new_AGEMA_signal_24404 ;
    wire new_AGEMA_signal_24405 ;
    wire new_AGEMA_signal_24406 ;
    wire new_AGEMA_signal_24407 ;
    wire new_AGEMA_signal_24408 ;
    wire new_AGEMA_signal_24409 ;
    wire new_AGEMA_signal_24410 ;
    wire new_AGEMA_signal_24411 ;
    wire new_AGEMA_signal_24412 ;
    wire new_AGEMA_signal_24413 ;
    wire new_AGEMA_signal_24414 ;
    wire new_AGEMA_signal_24415 ;
    wire new_AGEMA_signal_24416 ;
    wire new_AGEMA_signal_24417 ;
    wire new_AGEMA_signal_24418 ;
    wire new_AGEMA_signal_24419 ;
    wire new_AGEMA_signal_24420 ;
    wire new_AGEMA_signal_24421 ;
    wire new_AGEMA_signal_24422 ;
    wire new_AGEMA_signal_24423 ;
    wire new_AGEMA_signal_24424 ;
    wire new_AGEMA_signal_24425 ;
    wire new_AGEMA_signal_24426 ;
    wire new_AGEMA_signal_24427 ;
    wire new_AGEMA_signal_24428 ;
    wire new_AGEMA_signal_24429 ;
    wire new_AGEMA_signal_24430 ;
    wire new_AGEMA_signal_24431 ;
    wire new_AGEMA_signal_24432 ;
    wire new_AGEMA_signal_24433 ;
    wire new_AGEMA_signal_24434 ;
    wire new_AGEMA_signal_24435 ;
    wire new_AGEMA_signal_24436 ;
    wire new_AGEMA_signal_24437 ;
    wire new_AGEMA_signal_24438 ;
    wire new_AGEMA_signal_24439 ;
    wire new_AGEMA_signal_24440 ;
    wire new_AGEMA_signal_24441 ;
    wire new_AGEMA_signal_24442 ;
    wire new_AGEMA_signal_24443 ;
    wire new_AGEMA_signal_24444 ;
    wire new_AGEMA_signal_24445 ;
    wire new_AGEMA_signal_24446 ;
    wire new_AGEMA_signal_24447 ;
    wire new_AGEMA_signal_24448 ;
    wire new_AGEMA_signal_24449 ;
    wire new_AGEMA_signal_24450 ;
    wire new_AGEMA_signal_24451 ;
    wire new_AGEMA_signal_24452 ;
    wire new_AGEMA_signal_24453 ;
    wire new_AGEMA_signal_24454 ;
    wire new_AGEMA_signal_24455 ;
    wire new_AGEMA_signal_24456 ;
    wire new_AGEMA_signal_24457 ;
    wire new_AGEMA_signal_24458 ;
    wire new_AGEMA_signal_24459 ;
    wire new_AGEMA_signal_24460 ;
    wire new_AGEMA_signal_24461 ;
    wire new_AGEMA_signal_24462 ;
    wire new_AGEMA_signal_24463 ;
    wire new_AGEMA_signal_24464 ;
    wire new_AGEMA_signal_24465 ;
    wire new_AGEMA_signal_24466 ;
    wire new_AGEMA_signal_24467 ;
    wire new_AGEMA_signal_24468 ;
    wire new_AGEMA_signal_24469 ;
    wire new_AGEMA_signal_24470 ;
    wire new_AGEMA_signal_24471 ;
    wire new_AGEMA_signal_24472 ;
    wire new_AGEMA_signal_24473 ;
    wire new_AGEMA_signal_24474 ;
    wire new_AGEMA_signal_24475 ;
    wire new_AGEMA_signal_24476 ;
    wire new_AGEMA_signal_24477 ;
    wire new_AGEMA_signal_24478 ;
    wire new_AGEMA_signal_24479 ;
    wire new_AGEMA_signal_24480 ;
    wire new_AGEMA_signal_24481 ;
    wire new_AGEMA_signal_24482 ;
    wire new_AGEMA_signal_24483 ;
    wire new_AGEMA_signal_24484 ;
    wire new_AGEMA_signal_24485 ;
    wire new_AGEMA_signal_24486 ;
    wire new_AGEMA_signal_24487 ;
    wire new_AGEMA_signal_24488 ;
    wire new_AGEMA_signal_24489 ;
    wire new_AGEMA_signal_24490 ;
    wire new_AGEMA_signal_24491 ;
    wire new_AGEMA_signal_24492 ;
    wire new_AGEMA_signal_24493 ;
    wire new_AGEMA_signal_24494 ;
    wire new_AGEMA_signal_24495 ;
    wire new_AGEMA_signal_24496 ;
    wire new_AGEMA_signal_24497 ;
    wire new_AGEMA_signal_24498 ;
    wire new_AGEMA_signal_24499 ;
    wire new_AGEMA_signal_24500 ;
    wire new_AGEMA_signal_24501 ;
    wire new_AGEMA_signal_24502 ;
    wire new_AGEMA_signal_24503 ;
    wire new_AGEMA_signal_24504 ;
    wire new_AGEMA_signal_24505 ;
    wire new_AGEMA_signal_24506 ;
    wire new_AGEMA_signal_24507 ;
    wire new_AGEMA_signal_24508 ;
    wire new_AGEMA_signal_24509 ;
    wire new_AGEMA_signal_24510 ;
    wire new_AGEMA_signal_24511 ;
    wire new_AGEMA_signal_24512 ;
    wire new_AGEMA_signal_24513 ;
    wire new_AGEMA_signal_24514 ;
    wire new_AGEMA_signal_24515 ;
    wire new_AGEMA_signal_24516 ;
    wire new_AGEMA_signal_24517 ;
    wire new_AGEMA_signal_24518 ;
    wire new_AGEMA_signal_24519 ;
    wire new_AGEMA_signal_24520 ;
    wire new_AGEMA_signal_24521 ;
    wire new_AGEMA_signal_24522 ;
    wire new_AGEMA_signal_24523 ;
    wire new_AGEMA_signal_24524 ;
    wire new_AGEMA_signal_24525 ;
    wire new_AGEMA_signal_24526 ;
    wire new_AGEMA_signal_24527 ;
    wire new_AGEMA_signal_24528 ;
    wire new_AGEMA_signal_24529 ;
    wire new_AGEMA_signal_24530 ;
    wire new_AGEMA_signal_24531 ;
    wire new_AGEMA_signal_24532 ;
    wire new_AGEMA_signal_24533 ;
    wire new_AGEMA_signal_24534 ;
    wire new_AGEMA_signal_24535 ;
    wire new_AGEMA_signal_24536 ;
    wire new_AGEMA_signal_24537 ;
    wire new_AGEMA_signal_24538 ;
    wire new_AGEMA_signal_24539 ;
    wire new_AGEMA_signal_24540 ;
    wire new_AGEMA_signal_24541 ;
    wire new_AGEMA_signal_24542 ;
    wire new_AGEMA_signal_24543 ;
    wire new_AGEMA_signal_24544 ;
    wire new_AGEMA_signal_24545 ;
    wire new_AGEMA_signal_24546 ;
    wire new_AGEMA_signal_24547 ;
    wire new_AGEMA_signal_24548 ;
    wire new_AGEMA_signal_24549 ;
    wire new_AGEMA_signal_24550 ;
    wire new_AGEMA_signal_24551 ;
    wire new_AGEMA_signal_24552 ;
    wire new_AGEMA_signal_24553 ;
    wire new_AGEMA_signal_24554 ;
    wire new_AGEMA_signal_24555 ;
    wire new_AGEMA_signal_24556 ;
    wire new_AGEMA_signal_24557 ;
    wire new_AGEMA_signal_24558 ;
    wire new_AGEMA_signal_24559 ;
    wire new_AGEMA_signal_24560 ;
    wire new_AGEMA_signal_24561 ;
    wire new_AGEMA_signal_24562 ;
    wire new_AGEMA_signal_24563 ;
    wire new_AGEMA_signal_24564 ;
    wire new_AGEMA_signal_24565 ;
    wire new_AGEMA_signal_24566 ;
    wire new_AGEMA_signal_24567 ;
    wire new_AGEMA_signal_24568 ;
    wire new_AGEMA_signal_24569 ;
    wire new_AGEMA_signal_24570 ;
    wire new_AGEMA_signal_24571 ;
    wire new_AGEMA_signal_24572 ;
    wire new_AGEMA_signal_24573 ;
    wire new_AGEMA_signal_24574 ;
    wire new_AGEMA_signal_24575 ;
    wire new_AGEMA_signal_24576 ;
    wire new_AGEMA_signal_24577 ;
    wire new_AGEMA_signal_24578 ;
    wire new_AGEMA_signal_24579 ;
    wire new_AGEMA_signal_24580 ;
    wire new_AGEMA_signal_24581 ;
    wire new_AGEMA_signal_24582 ;
    wire new_AGEMA_signal_24583 ;
    wire new_AGEMA_signal_24584 ;
    wire new_AGEMA_signal_24585 ;
    wire new_AGEMA_signal_24586 ;
    wire new_AGEMA_signal_24587 ;
    wire new_AGEMA_signal_24588 ;
    wire new_AGEMA_signal_24589 ;
    wire new_AGEMA_signal_24590 ;
    wire new_AGEMA_signal_24591 ;
    wire new_AGEMA_signal_24592 ;
    wire new_AGEMA_signal_24593 ;
    wire new_AGEMA_signal_24594 ;
    wire new_AGEMA_signal_24595 ;
    wire new_AGEMA_signal_24596 ;
    wire new_AGEMA_signal_24597 ;
    wire new_AGEMA_signal_24598 ;
    wire new_AGEMA_signal_24599 ;
    wire new_AGEMA_signal_24600 ;
    wire new_AGEMA_signal_24601 ;
    wire new_AGEMA_signal_24602 ;
    wire new_AGEMA_signal_24603 ;
    wire new_AGEMA_signal_24604 ;
    wire new_AGEMA_signal_24605 ;
    wire new_AGEMA_signal_24606 ;
    wire new_AGEMA_signal_24607 ;
    wire new_AGEMA_signal_24608 ;
    wire new_AGEMA_signal_24609 ;
    wire new_AGEMA_signal_24610 ;
    wire new_AGEMA_signal_24611 ;
    wire new_AGEMA_signal_24612 ;
    wire new_AGEMA_signal_24613 ;
    wire new_AGEMA_signal_24614 ;
    wire new_AGEMA_signal_24615 ;
    wire new_AGEMA_signal_24616 ;
    wire new_AGEMA_signal_24617 ;
    wire new_AGEMA_signal_24618 ;
    wire new_AGEMA_signal_24619 ;
    wire new_AGEMA_signal_24620 ;
    wire new_AGEMA_signal_24621 ;
    wire new_AGEMA_signal_24622 ;
    wire new_AGEMA_signal_24623 ;
    wire new_AGEMA_signal_24624 ;
    wire new_AGEMA_signal_24625 ;
    wire new_AGEMA_signal_24626 ;
    wire new_AGEMA_signal_24627 ;
    wire new_AGEMA_signal_24628 ;
    wire new_AGEMA_signal_24629 ;
    wire new_AGEMA_signal_24630 ;
    wire new_AGEMA_signal_24631 ;
    wire new_AGEMA_signal_24632 ;
    wire new_AGEMA_signal_24633 ;
    wire new_AGEMA_signal_24634 ;
    wire new_AGEMA_signal_24635 ;
    wire new_AGEMA_signal_24636 ;
    wire new_AGEMA_signal_24637 ;
    wire new_AGEMA_signal_24638 ;
    wire new_AGEMA_signal_24639 ;
    wire new_AGEMA_signal_24640 ;
    wire new_AGEMA_signal_24641 ;
    wire new_AGEMA_signal_24642 ;
    wire new_AGEMA_signal_24643 ;
    wire new_AGEMA_signal_24644 ;
    wire new_AGEMA_signal_24645 ;
    wire new_AGEMA_signal_24646 ;
    wire new_AGEMA_signal_24647 ;
    wire new_AGEMA_signal_24648 ;
    wire new_AGEMA_signal_24649 ;
    wire new_AGEMA_signal_24650 ;
    wire new_AGEMA_signal_24651 ;
    wire new_AGEMA_signal_24652 ;
    wire new_AGEMA_signal_24653 ;
    wire new_AGEMA_signal_24654 ;
    wire new_AGEMA_signal_24655 ;
    wire new_AGEMA_signal_24656 ;
    wire new_AGEMA_signal_24657 ;
    wire new_AGEMA_signal_24658 ;
    wire new_AGEMA_signal_24659 ;
    wire new_AGEMA_signal_24660 ;
    wire new_AGEMA_signal_24661 ;
    wire new_AGEMA_signal_24662 ;
    wire new_AGEMA_signal_24663 ;
    wire new_AGEMA_signal_24664 ;
    wire new_AGEMA_signal_24665 ;
    wire new_AGEMA_signal_24666 ;
    wire new_AGEMA_signal_24667 ;
    wire new_AGEMA_signal_24668 ;
    wire new_AGEMA_signal_24669 ;
    wire new_AGEMA_signal_24670 ;
    wire new_AGEMA_signal_24671 ;
    wire new_AGEMA_signal_24672 ;
    wire new_AGEMA_signal_24673 ;
    wire new_AGEMA_signal_24674 ;
    wire new_AGEMA_signal_24675 ;
    wire new_AGEMA_signal_24676 ;
    wire new_AGEMA_signal_24677 ;
    wire new_AGEMA_signal_24678 ;
    wire new_AGEMA_signal_24679 ;
    wire new_AGEMA_signal_24680 ;
    wire new_AGEMA_signal_24681 ;
    wire new_AGEMA_signal_24682 ;
    wire new_AGEMA_signal_24683 ;
    wire new_AGEMA_signal_24684 ;
    wire new_AGEMA_signal_24685 ;
    wire new_AGEMA_signal_24686 ;
    wire new_AGEMA_signal_24687 ;
    wire new_AGEMA_signal_24688 ;
    wire new_AGEMA_signal_24689 ;
    wire new_AGEMA_signal_24690 ;
    wire new_AGEMA_signal_24691 ;
    wire new_AGEMA_signal_24692 ;
    wire new_AGEMA_signal_24693 ;
    wire new_AGEMA_signal_24694 ;
    wire new_AGEMA_signal_24695 ;
    wire new_AGEMA_signal_24696 ;
    wire new_AGEMA_signal_24697 ;
    wire new_AGEMA_signal_24698 ;
    wire new_AGEMA_signal_24699 ;
    wire new_AGEMA_signal_24700 ;
    wire new_AGEMA_signal_24701 ;
    wire new_AGEMA_signal_24702 ;
    wire new_AGEMA_signal_24703 ;
    wire new_AGEMA_signal_24704 ;
    wire new_AGEMA_signal_24705 ;
    wire new_AGEMA_signal_24706 ;
    wire new_AGEMA_signal_24707 ;
    wire new_AGEMA_signal_24708 ;
    wire new_AGEMA_signal_24709 ;
    wire new_AGEMA_signal_24710 ;
    wire new_AGEMA_signal_24711 ;
    wire new_AGEMA_signal_24712 ;
    wire new_AGEMA_signal_24713 ;
    wire new_AGEMA_signal_24714 ;
    wire new_AGEMA_signal_24715 ;
    wire new_AGEMA_signal_24716 ;
    wire new_AGEMA_signal_24717 ;
    wire new_AGEMA_signal_24718 ;
    wire new_AGEMA_signal_24719 ;
    wire new_AGEMA_signal_24720 ;
    wire new_AGEMA_signal_24721 ;
    wire new_AGEMA_signal_24722 ;
    wire new_AGEMA_signal_24723 ;
    wire new_AGEMA_signal_24724 ;
    wire new_AGEMA_signal_24725 ;
    wire new_AGEMA_signal_24726 ;
    wire new_AGEMA_signal_24727 ;
    wire new_AGEMA_signal_24728 ;
    wire new_AGEMA_signal_24729 ;
    wire new_AGEMA_signal_24730 ;
    wire new_AGEMA_signal_24731 ;
    wire new_AGEMA_signal_24732 ;
    wire new_AGEMA_signal_24733 ;
    wire new_AGEMA_signal_24734 ;
    wire new_AGEMA_signal_24735 ;
    wire new_AGEMA_signal_24736 ;
    wire new_AGEMA_signal_24737 ;
    wire new_AGEMA_signal_24738 ;
    wire new_AGEMA_signal_24739 ;
    wire new_AGEMA_signal_24740 ;
    wire new_AGEMA_signal_24741 ;
    wire new_AGEMA_signal_24742 ;
    wire new_AGEMA_signal_24743 ;
    wire new_AGEMA_signal_24744 ;
    wire new_AGEMA_signal_24745 ;
    wire new_AGEMA_signal_24746 ;
    wire new_AGEMA_signal_24747 ;
    wire new_AGEMA_signal_24748 ;
    wire new_AGEMA_signal_24749 ;
    wire new_AGEMA_signal_24750 ;
    wire new_AGEMA_signal_24751 ;
    wire new_AGEMA_signal_24752 ;
    wire new_AGEMA_signal_24753 ;
    wire new_AGEMA_signal_24754 ;
    wire new_AGEMA_signal_24755 ;
    wire new_AGEMA_signal_24756 ;
    wire new_AGEMA_signal_24757 ;
    wire new_AGEMA_signal_24758 ;
    wire new_AGEMA_signal_24759 ;
    wire new_AGEMA_signal_24760 ;
    wire new_AGEMA_signal_24761 ;
    wire new_AGEMA_signal_24762 ;
    wire new_AGEMA_signal_24763 ;
    wire new_AGEMA_signal_24764 ;
    wire new_AGEMA_signal_24765 ;
    wire new_AGEMA_signal_24766 ;
    wire new_AGEMA_signal_24767 ;
    wire new_AGEMA_signal_24768 ;
    wire new_AGEMA_signal_24769 ;
    wire new_AGEMA_signal_24770 ;
    wire new_AGEMA_signal_24771 ;
    wire new_AGEMA_signal_24772 ;
    wire new_AGEMA_signal_24773 ;
    wire new_AGEMA_signal_24774 ;
    wire new_AGEMA_signal_24775 ;
    wire new_AGEMA_signal_24776 ;
    wire new_AGEMA_signal_24777 ;
    wire new_AGEMA_signal_24778 ;
    wire new_AGEMA_signal_24779 ;
    wire new_AGEMA_signal_24780 ;
    wire new_AGEMA_signal_24781 ;
    wire new_AGEMA_signal_24782 ;
    wire new_AGEMA_signal_24783 ;
    wire new_AGEMA_signal_24784 ;
    wire new_AGEMA_signal_24785 ;
    wire new_AGEMA_signal_24786 ;
    wire new_AGEMA_signal_24787 ;
    wire new_AGEMA_signal_24788 ;
    wire new_AGEMA_signal_24789 ;
    wire new_AGEMA_signal_24790 ;
    wire new_AGEMA_signal_24791 ;
    wire new_AGEMA_signal_24792 ;
    wire new_AGEMA_signal_24793 ;
    wire new_AGEMA_signal_24794 ;
    wire new_AGEMA_signal_24795 ;
    wire new_AGEMA_signal_24796 ;
    wire new_AGEMA_signal_24797 ;
    wire new_AGEMA_signal_24798 ;
    wire new_AGEMA_signal_24799 ;
    wire new_AGEMA_signal_24800 ;
    wire new_AGEMA_signal_24801 ;
    wire new_AGEMA_signal_24802 ;
    wire new_AGEMA_signal_24803 ;
    wire new_AGEMA_signal_24804 ;
    wire new_AGEMA_signal_24805 ;
    wire new_AGEMA_signal_24806 ;
    wire new_AGEMA_signal_24807 ;
    wire new_AGEMA_signal_24808 ;
    wire new_AGEMA_signal_24809 ;
    wire new_AGEMA_signal_24810 ;
    wire new_AGEMA_signal_24811 ;
    wire new_AGEMA_signal_24812 ;
    wire new_AGEMA_signal_24813 ;
    wire new_AGEMA_signal_24814 ;
    wire new_AGEMA_signal_24815 ;
    wire new_AGEMA_signal_24816 ;
    wire new_AGEMA_signal_24817 ;
    wire new_AGEMA_signal_24818 ;
    wire new_AGEMA_signal_24819 ;
    wire new_AGEMA_signal_24820 ;
    wire new_AGEMA_signal_24821 ;
    wire new_AGEMA_signal_24822 ;
    wire new_AGEMA_signal_24823 ;
    wire new_AGEMA_signal_24824 ;
    wire new_AGEMA_signal_24825 ;
    wire new_AGEMA_signal_24826 ;
    wire new_AGEMA_signal_24827 ;
    wire new_AGEMA_signal_24828 ;
    wire new_AGEMA_signal_24829 ;
    wire new_AGEMA_signal_24830 ;
    wire new_AGEMA_signal_24831 ;
    wire new_AGEMA_signal_24832 ;
    wire new_AGEMA_signal_24833 ;
    wire new_AGEMA_signal_24834 ;
    wire new_AGEMA_signal_24835 ;
    wire new_AGEMA_signal_24836 ;
    wire new_AGEMA_signal_24837 ;
    wire new_AGEMA_signal_24838 ;
    wire new_AGEMA_signal_24839 ;
    wire new_AGEMA_signal_24840 ;
    wire new_AGEMA_signal_24841 ;
    wire new_AGEMA_signal_24842 ;
    wire new_AGEMA_signal_24843 ;
    wire new_AGEMA_signal_24844 ;
    wire new_AGEMA_signal_24845 ;
    wire new_AGEMA_signal_24846 ;
    wire new_AGEMA_signal_24847 ;
    wire new_AGEMA_signal_24848 ;
    wire new_AGEMA_signal_24849 ;
    wire new_AGEMA_signal_24850 ;
    wire new_AGEMA_signal_24851 ;
    wire new_AGEMA_signal_24852 ;
    wire new_AGEMA_signal_24853 ;
    wire new_AGEMA_signal_24854 ;
    wire new_AGEMA_signal_24855 ;
    wire new_AGEMA_signal_24856 ;
    wire new_AGEMA_signal_24857 ;
    wire new_AGEMA_signal_24858 ;
    wire new_AGEMA_signal_24859 ;
    wire new_AGEMA_signal_24860 ;
    wire new_AGEMA_signal_24861 ;
    wire new_AGEMA_signal_24862 ;
    wire new_AGEMA_signal_24863 ;
    wire new_AGEMA_signal_24864 ;
    wire new_AGEMA_signal_24865 ;
    wire new_AGEMA_signal_24866 ;
    wire new_AGEMA_signal_24867 ;
    wire new_AGEMA_signal_24868 ;
    wire new_AGEMA_signal_24869 ;
    wire new_AGEMA_signal_24870 ;
    wire new_AGEMA_signal_24871 ;
    wire new_AGEMA_signal_24872 ;
    wire new_AGEMA_signal_24873 ;
    wire new_AGEMA_signal_24874 ;
    wire new_AGEMA_signal_24875 ;
    wire new_AGEMA_signal_24876 ;
    wire new_AGEMA_signal_24877 ;
    wire new_AGEMA_signal_24878 ;
    wire new_AGEMA_signal_24879 ;
    wire new_AGEMA_signal_24880 ;
    wire new_AGEMA_signal_24881 ;
    wire new_AGEMA_signal_24882 ;
    wire new_AGEMA_signal_24883 ;
    wire new_AGEMA_signal_24884 ;
    wire new_AGEMA_signal_24885 ;
    wire new_AGEMA_signal_24886 ;
    wire new_AGEMA_signal_24887 ;
    wire new_AGEMA_signal_24888 ;
    wire new_AGEMA_signal_24889 ;
    wire new_AGEMA_signal_24890 ;
    wire new_AGEMA_signal_24891 ;
    wire new_AGEMA_signal_24892 ;
    wire new_AGEMA_signal_24893 ;
    wire new_AGEMA_signal_24894 ;
    wire new_AGEMA_signal_24895 ;
    wire new_AGEMA_signal_24896 ;
    wire new_AGEMA_signal_24897 ;
    wire new_AGEMA_signal_24898 ;
    wire new_AGEMA_signal_24899 ;
    wire new_AGEMA_signal_24900 ;
    wire new_AGEMA_signal_24901 ;
    wire new_AGEMA_signal_24902 ;
    wire new_AGEMA_signal_24903 ;
    wire new_AGEMA_signal_24904 ;
    wire new_AGEMA_signal_24905 ;
    wire new_AGEMA_signal_24906 ;
    wire new_AGEMA_signal_24907 ;
    wire new_AGEMA_signal_24908 ;
    wire new_AGEMA_signal_24909 ;
    wire new_AGEMA_signal_24910 ;
    wire new_AGEMA_signal_24911 ;
    wire new_AGEMA_signal_24912 ;
    wire new_AGEMA_signal_24913 ;
    wire new_AGEMA_signal_24914 ;
    wire new_AGEMA_signal_24915 ;
    wire new_AGEMA_signal_24916 ;
    wire new_AGEMA_signal_24917 ;
    wire new_AGEMA_signal_24918 ;
    wire new_AGEMA_signal_24919 ;
    wire new_AGEMA_signal_24920 ;
    wire new_AGEMA_signal_24921 ;
    wire new_AGEMA_signal_24922 ;
    wire new_AGEMA_signal_24923 ;
    wire new_AGEMA_signal_24924 ;
    wire new_AGEMA_signal_24925 ;
    wire new_AGEMA_signal_24926 ;
    wire new_AGEMA_signal_24927 ;
    wire new_AGEMA_signal_24928 ;
    wire new_AGEMA_signal_24929 ;
    wire new_AGEMA_signal_24930 ;
    wire new_AGEMA_signal_24931 ;
    wire new_AGEMA_signal_24932 ;
    wire new_AGEMA_signal_24933 ;
    wire new_AGEMA_signal_24934 ;
    wire new_AGEMA_signal_24935 ;
    wire new_AGEMA_signal_24936 ;
    wire new_AGEMA_signal_24937 ;
    wire new_AGEMA_signal_24938 ;
    wire new_AGEMA_signal_24939 ;
    wire new_AGEMA_signal_24940 ;
    wire new_AGEMA_signal_24941 ;
    wire new_AGEMA_signal_24942 ;
    wire new_AGEMA_signal_24943 ;
    wire new_AGEMA_signal_24944 ;
    wire new_AGEMA_signal_24945 ;
    wire new_AGEMA_signal_24946 ;
    wire new_AGEMA_signal_24947 ;
    wire new_AGEMA_signal_24948 ;
    wire new_AGEMA_signal_24949 ;
    wire new_AGEMA_signal_24950 ;
    wire new_AGEMA_signal_24951 ;
    wire new_AGEMA_signal_24952 ;
    wire new_AGEMA_signal_24953 ;
    wire new_AGEMA_signal_24954 ;
    wire new_AGEMA_signal_24955 ;
    wire new_AGEMA_signal_24956 ;
    wire new_AGEMA_signal_24957 ;
    wire new_AGEMA_signal_24958 ;
    wire new_AGEMA_signal_24959 ;
    wire new_AGEMA_signal_24960 ;
    wire new_AGEMA_signal_24961 ;
    wire new_AGEMA_signal_24962 ;
    wire new_AGEMA_signal_24963 ;
    wire new_AGEMA_signal_24964 ;
    wire new_AGEMA_signal_24965 ;
    wire new_AGEMA_signal_24966 ;
    wire new_AGEMA_signal_24967 ;
    wire new_AGEMA_signal_24968 ;
    wire new_AGEMA_signal_24969 ;
    wire new_AGEMA_signal_24970 ;
    wire new_AGEMA_signal_24971 ;
    wire new_AGEMA_signal_24972 ;
    wire new_AGEMA_signal_24973 ;
    wire new_AGEMA_signal_24974 ;
    wire new_AGEMA_signal_24975 ;
    wire new_AGEMA_signal_24976 ;
    wire new_AGEMA_signal_24977 ;
    wire new_AGEMA_signal_24978 ;
    wire new_AGEMA_signal_24979 ;
    wire new_AGEMA_signal_24980 ;
    wire new_AGEMA_signal_24981 ;
    wire new_AGEMA_signal_24982 ;
    wire new_AGEMA_signal_24983 ;
    wire new_AGEMA_signal_24984 ;
    wire new_AGEMA_signal_24985 ;
    wire new_AGEMA_signal_24986 ;
    wire new_AGEMA_signal_24987 ;
    wire new_AGEMA_signal_24988 ;
    wire new_AGEMA_signal_24989 ;
    wire new_AGEMA_signal_24990 ;
    wire new_AGEMA_signal_24991 ;
    wire new_AGEMA_signal_24992 ;
    wire new_AGEMA_signal_24993 ;
    wire new_AGEMA_signal_24994 ;
    wire new_AGEMA_signal_24995 ;
    wire new_AGEMA_signal_24996 ;
    wire new_AGEMA_signal_24997 ;
    wire new_AGEMA_signal_24998 ;
    wire new_AGEMA_signal_24999 ;
    wire new_AGEMA_signal_25000 ;
    wire new_AGEMA_signal_25001 ;
    wire new_AGEMA_signal_25002 ;
    wire new_AGEMA_signal_25003 ;
    wire new_AGEMA_signal_25004 ;
    wire new_AGEMA_signal_25005 ;
    wire new_AGEMA_signal_25006 ;
    wire new_AGEMA_signal_25007 ;
    wire new_AGEMA_signal_25008 ;
    wire new_AGEMA_signal_25009 ;
    wire new_AGEMA_signal_25010 ;
    wire new_AGEMA_signal_25011 ;
    wire new_AGEMA_signal_25012 ;
    wire new_AGEMA_signal_25013 ;
    wire new_AGEMA_signal_25014 ;
    wire new_AGEMA_signal_25015 ;
    wire new_AGEMA_signal_25016 ;
    wire new_AGEMA_signal_25017 ;
    wire new_AGEMA_signal_25018 ;
    wire new_AGEMA_signal_25019 ;
    wire new_AGEMA_signal_25020 ;
    wire new_AGEMA_signal_25021 ;
    wire new_AGEMA_signal_25022 ;
    wire new_AGEMA_signal_25023 ;
    wire new_AGEMA_signal_25024 ;
    wire new_AGEMA_signal_25025 ;
    wire new_AGEMA_signal_25026 ;
    wire new_AGEMA_signal_25027 ;
    wire new_AGEMA_signal_25028 ;
    wire new_AGEMA_signal_25029 ;
    wire new_AGEMA_signal_25030 ;
    wire new_AGEMA_signal_25031 ;
    wire new_AGEMA_signal_25032 ;
    wire new_AGEMA_signal_25033 ;
    wire new_AGEMA_signal_25034 ;
    wire new_AGEMA_signal_25035 ;
    wire new_AGEMA_signal_25036 ;
    wire new_AGEMA_signal_25037 ;
    wire new_AGEMA_signal_25038 ;
    wire new_AGEMA_signal_25039 ;
    wire new_AGEMA_signal_25040 ;
    wire new_AGEMA_signal_25041 ;
    wire new_AGEMA_signal_25042 ;
    wire new_AGEMA_signal_25043 ;
    wire new_AGEMA_signal_25044 ;
    wire new_AGEMA_signal_25045 ;
    wire new_AGEMA_signal_25046 ;
    wire new_AGEMA_signal_25047 ;
    wire new_AGEMA_signal_25048 ;
    wire new_AGEMA_signal_25049 ;
    wire new_AGEMA_signal_25050 ;
    wire new_AGEMA_signal_25051 ;
    wire new_AGEMA_signal_25052 ;
    wire new_AGEMA_signal_25053 ;
    wire new_AGEMA_signal_25054 ;
    wire new_AGEMA_signal_25055 ;
    wire new_AGEMA_signal_25056 ;
    wire new_AGEMA_signal_25057 ;
    wire new_AGEMA_signal_25058 ;
    wire new_AGEMA_signal_25059 ;
    wire new_AGEMA_signal_25060 ;
    wire new_AGEMA_signal_25061 ;
    wire new_AGEMA_signal_25062 ;
    wire new_AGEMA_signal_25063 ;
    wire new_AGEMA_signal_25064 ;
    wire new_AGEMA_signal_25065 ;
    wire new_AGEMA_signal_25066 ;
    wire new_AGEMA_signal_25067 ;
    wire new_AGEMA_signal_25068 ;
    wire new_AGEMA_signal_25069 ;
    wire new_AGEMA_signal_25070 ;
    wire new_AGEMA_signal_25071 ;
    wire new_AGEMA_signal_25072 ;
    wire new_AGEMA_signal_25073 ;
    wire new_AGEMA_signal_25074 ;
    wire new_AGEMA_signal_25075 ;
    wire new_AGEMA_signal_25076 ;
    wire new_AGEMA_signal_25077 ;
    wire new_AGEMA_signal_25078 ;
    wire new_AGEMA_signal_25079 ;
    wire new_AGEMA_signal_25080 ;
    wire new_AGEMA_signal_25081 ;
    wire new_AGEMA_signal_25082 ;
    wire new_AGEMA_signal_25083 ;
    wire new_AGEMA_signal_25084 ;
    wire new_AGEMA_signal_25085 ;
    wire new_AGEMA_signal_25086 ;
    wire new_AGEMA_signal_25087 ;
    wire new_AGEMA_signal_25088 ;
    wire new_AGEMA_signal_25089 ;
    wire new_AGEMA_signal_25090 ;
    wire new_AGEMA_signal_25091 ;
    wire new_AGEMA_signal_25092 ;
    wire new_AGEMA_signal_25093 ;
    wire new_AGEMA_signal_25094 ;
    wire new_AGEMA_signal_25095 ;
    wire new_AGEMA_signal_25096 ;
    wire new_AGEMA_signal_25097 ;
    wire new_AGEMA_signal_25098 ;
    wire new_AGEMA_signal_25099 ;
    wire new_AGEMA_signal_25100 ;
    wire new_AGEMA_signal_25101 ;
    wire new_AGEMA_signal_25102 ;
    wire new_AGEMA_signal_25103 ;
    wire new_AGEMA_signal_25104 ;
    wire new_AGEMA_signal_25105 ;
    wire new_AGEMA_signal_25106 ;
    wire new_AGEMA_signal_25107 ;
    wire new_AGEMA_signal_25108 ;
    wire new_AGEMA_signal_25109 ;
    wire new_AGEMA_signal_25110 ;
    wire new_AGEMA_signal_25111 ;
    wire new_AGEMA_signal_25112 ;
    wire new_AGEMA_signal_25113 ;
    wire new_AGEMA_signal_25114 ;
    wire new_AGEMA_signal_25115 ;
    wire new_AGEMA_signal_25116 ;
    wire new_AGEMA_signal_25117 ;
    wire new_AGEMA_signal_25118 ;
    wire new_AGEMA_signal_25119 ;
    wire new_AGEMA_signal_25120 ;
    wire new_AGEMA_signal_25121 ;
    wire new_AGEMA_signal_25122 ;
    wire new_AGEMA_signal_25123 ;
    wire new_AGEMA_signal_25124 ;
    wire new_AGEMA_signal_25125 ;
    wire new_AGEMA_signal_25126 ;
    wire new_AGEMA_signal_25127 ;
    wire new_AGEMA_signal_25128 ;
    wire new_AGEMA_signal_25129 ;
    wire new_AGEMA_signal_25130 ;
    wire new_AGEMA_signal_25131 ;
    wire new_AGEMA_signal_25132 ;
    wire new_AGEMA_signal_25133 ;
    wire new_AGEMA_signal_25134 ;
    wire new_AGEMA_signal_25135 ;
    wire new_AGEMA_signal_25136 ;
    wire new_AGEMA_signal_25137 ;
    wire new_AGEMA_signal_25138 ;
    wire new_AGEMA_signal_25139 ;
    wire new_AGEMA_signal_25140 ;
    wire new_AGEMA_signal_25141 ;
    wire new_AGEMA_signal_25142 ;
    wire new_AGEMA_signal_25143 ;
    wire new_AGEMA_signal_25144 ;
    wire new_AGEMA_signal_25145 ;
    wire new_AGEMA_signal_25146 ;
    wire new_AGEMA_signal_25147 ;
    wire new_AGEMA_signal_25148 ;
    wire new_AGEMA_signal_25149 ;
    wire new_AGEMA_signal_25150 ;
    wire new_AGEMA_signal_25151 ;
    wire new_AGEMA_signal_25152 ;
    wire new_AGEMA_signal_25153 ;
    wire new_AGEMA_signal_25154 ;
    wire new_AGEMA_signal_25155 ;
    wire new_AGEMA_signal_25156 ;
    wire new_AGEMA_signal_25157 ;
    wire new_AGEMA_signal_25158 ;
    wire new_AGEMA_signal_25159 ;
    wire new_AGEMA_signal_25160 ;
    wire new_AGEMA_signal_25161 ;
    wire new_AGEMA_signal_25162 ;
    wire new_AGEMA_signal_25163 ;
    wire new_AGEMA_signal_25164 ;
    wire new_AGEMA_signal_25165 ;
    wire new_AGEMA_signal_25166 ;
    wire new_AGEMA_signal_25167 ;
    wire new_AGEMA_signal_25168 ;
    wire new_AGEMA_signal_25169 ;
    wire new_AGEMA_signal_25170 ;
    wire new_AGEMA_signal_25171 ;
    wire new_AGEMA_signal_25172 ;
    wire new_AGEMA_signal_25173 ;
    wire new_AGEMA_signal_25174 ;
    wire new_AGEMA_signal_25175 ;
    wire new_AGEMA_signal_25176 ;
    wire new_AGEMA_signal_25177 ;
    wire new_AGEMA_signal_25178 ;
    wire new_AGEMA_signal_25179 ;
    wire new_AGEMA_signal_25180 ;
    wire new_AGEMA_signal_25181 ;
    wire new_AGEMA_signal_25182 ;
    wire new_AGEMA_signal_25183 ;
    wire new_AGEMA_signal_25184 ;
    wire new_AGEMA_signal_25185 ;
    wire new_AGEMA_signal_25186 ;
    wire new_AGEMA_signal_25187 ;
    wire new_AGEMA_signal_25188 ;
    wire new_AGEMA_signal_25189 ;
    wire new_AGEMA_signal_25190 ;
    wire new_AGEMA_signal_25191 ;
    wire new_AGEMA_signal_25192 ;
    wire new_AGEMA_signal_25193 ;
    wire new_AGEMA_signal_25194 ;
    wire new_AGEMA_signal_25195 ;
    wire new_AGEMA_signal_25196 ;
    wire new_AGEMA_signal_25197 ;
    wire new_AGEMA_signal_25198 ;
    wire new_AGEMA_signal_25199 ;
    wire new_AGEMA_signal_25200 ;
    wire new_AGEMA_signal_25201 ;
    wire new_AGEMA_signal_25202 ;
    wire new_AGEMA_signal_25203 ;
    wire new_AGEMA_signal_25204 ;
    wire new_AGEMA_signal_25205 ;
    wire new_AGEMA_signal_25206 ;
    wire new_AGEMA_signal_25207 ;
    wire new_AGEMA_signal_25208 ;
    wire new_AGEMA_signal_25209 ;
    wire new_AGEMA_signal_25210 ;
    wire new_AGEMA_signal_25211 ;
    wire new_AGEMA_signal_25212 ;
    wire new_AGEMA_signal_25213 ;
    wire new_AGEMA_signal_25214 ;
    wire new_AGEMA_signal_25215 ;
    wire new_AGEMA_signal_25216 ;
    wire new_AGEMA_signal_25217 ;
    wire new_AGEMA_signal_25218 ;
    wire new_AGEMA_signal_25219 ;
    wire new_AGEMA_signal_25220 ;
    wire new_AGEMA_signal_25221 ;
    wire new_AGEMA_signal_25222 ;
    wire new_AGEMA_signal_25223 ;
    wire new_AGEMA_signal_25224 ;
    wire new_AGEMA_signal_25225 ;
    wire new_AGEMA_signal_25226 ;
    wire new_AGEMA_signal_25227 ;
    wire new_AGEMA_signal_25228 ;
    wire new_AGEMA_signal_25229 ;
    wire new_AGEMA_signal_25230 ;
    wire new_AGEMA_signal_25231 ;
    wire new_AGEMA_signal_25232 ;
    wire new_AGEMA_signal_25233 ;
    wire new_AGEMA_signal_25234 ;
    wire new_AGEMA_signal_25235 ;
    wire new_AGEMA_signal_25236 ;
    wire new_AGEMA_signal_25237 ;
    wire new_AGEMA_signal_25238 ;
    wire new_AGEMA_signal_25239 ;
    wire new_AGEMA_signal_25240 ;
    wire new_AGEMA_signal_25241 ;
    wire new_AGEMA_signal_25242 ;
    wire new_AGEMA_signal_25243 ;
    wire new_AGEMA_signal_25244 ;
    wire new_AGEMA_signal_25245 ;
    wire new_AGEMA_signal_25246 ;
    wire new_AGEMA_signal_25247 ;
    wire new_AGEMA_signal_25248 ;
    wire new_AGEMA_signal_25249 ;
    wire new_AGEMA_signal_25250 ;
    wire new_AGEMA_signal_25251 ;
    wire new_AGEMA_signal_25252 ;
    wire new_AGEMA_signal_25253 ;
    wire new_AGEMA_signal_25254 ;
    wire new_AGEMA_signal_25255 ;
    wire new_AGEMA_signal_25256 ;
    wire new_AGEMA_signal_25257 ;
    wire new_AGEMA_signal_25258 ;
    wire new_AGEMA_signal_25259 ;
    wire new_AGEMA_signal_25260 ;
    wire new_AGEMA_signal_25261 ;
    wire new_AGEMA_signal_25262 ;
    wire new_AGEMA_signal_25263 ;
    wire new_AGEMA_signal_25264 ;
    wire new_AGEMA_signal_25265 ;
    wire new_AGEMA_signal_25266 ;
    wire new_AGEMA_signal_25267 ;
    wire new_AGEMA_signal_25268 ;
    wire new_AGEMA_signal_25269 ;
    wire new_AGEMA_signal_25270 ;
    wire new_AGEMA_signal_25271 ;
    wire new_AGEMA_signal_25272 ;
    wire new_AGEMA_signal_25273 ;
    wire new_AGEMA_signal_25274 ;
    wire new_AGEMA_signal_25275 ;
    wire new_AGEMA_signal_25276 ;
    wire new_AGEMA_signal_25277 ;
    wire new_AGEMA_signal_25278 ;
    wire new_AGEMA_signal_25279 ;
    wire new_AGEMA_signal_25280 ;
    wire new_AGEMA_signal_25281 ;
    wire new_AGEMA_signal_25282 ;
    wire new_AGEMA_signal_25283 ;
    wire new_AGEMA_signal_25284 ;
    wire new_AGEMA_signal_25285 ;
    wire new_AGEMA_signal_25286 ;
    wire new_AGEMA_signal_25287 ;
    wire new_AGEMA_signal_25288 ;
    wire new_AGEMA_signal_25289 ;
    wire new_AGEMA_signal_25290 ;
    wire new_AGEMA_signal_25291 ;
    wire new_AGEMA_signal_25292 ;
    wire new_AGEMA_signal_25293 ;
    wire new_AGEMA_signal_25294 ;
    wire new_AGEMA_signal_25295 ;
    wire new_AGEMA_signal_25296 ;
    wire new_AGEMA_signal_25297 ;
    wire new_AGEMA_signal_25298 ;
    wire new_AGEMA_signal_25299 ;
    wire new_AGEMA_signal_25300 ;
    wire new_AGEMA_signal_25301 ;
    wire new_AGEMA_signal_25302 ;
    wire new_AGEMA_signal_25303 ;
    wire new_AGEMA_signal_25304 ;
    wire new_AGEMA_signal_25305 ;
    wire new_AGEMA_signal_25306 ;
    wire new_AGEMA_signal_25307 ;
    wire new_AGEMA_signal_25308 ;
    wire new_AGEMA_signal_25309 ;
    wire new_AGEMA_signal_25310 ;
    wire new_AGEMA_signal_25311 ;
    wire new_AGEMA_signal_25312 ;
    wire new_AGEMA_signal_25313 ;
    wire new_AGEMA_signal_25314 ;
    wire new_AGEMA_signal_25315 ;
    wire new_AGEMA_signal_25316 ;
    wire new_AGEMA_signal_25317 ;
    wire new_AGEMA_signal_25318 ;
    wire new_AGEMA_signal_25319 ;
    wire new_AGEMA_signal_25320 ;
    wire new_AGEMA_signal_25321 ;
    wire new_AGEMA_signal_25322 ;
    wire new_AGEMA_signal_25323 ;
    wire new_AGEMA_signal_25324 ;
    wire new_AGEMA_signal_25325 ;
    wire new_AGEMA_signal_25326 ;
    wire new_AGEMA_signal_25327 ;
    wire new_AGEMA_signal_25328 ;
    wire new_AGEMA_signal_25329 ;
    wire new_AGEMA_signal_25330 ;
    wire new_AGEMA_signal_25331 ;
    wire new_AGEMA_signal_25332 ;
    wire new_AGEMA_signal_25333 ;
    wire new_AGEMA_signal_25334 ;
    wire new_AGEMA_signal_25335 ;
    wire new_AGEMA_signal_25336 ;
    wire new_AGEMA_signal_25337 ;
    wire new_AGEMA_signal_25338 ;
    wire new_AGEMA_signal_25339 ;
    wire new_AGEMA_signal_25340 ;
    wire new_AGEMA_signal_25341 ;
    wire new_AGEMA_signal_25342 ;
    wire new_AGEMA_signal_25343 ;
    wire new_AGEMA_signal_25344 ;
    wire new_AGEMA_signal_25345 ;
    wire new_AGEMA_signal_25346 ;
    wire new_AGEMA_signal_25347 ;
    wire new_AGEMA_signal_25348 ;
    wire new_AGEMA_signal_25349 ;
    wire new_AGEMA_signal_25350 ;
    wire new_AGEMA_signal_25351 ;
    wire new_AGEMA_signal_25352 ;
    wire new_AGEMA_signal_25353 ;
    wire new_AGEMA_signal_25354 ;
    wire new_AGEMA_signal_25355 ;
    wire new_AGEMA_signal_25356 ;
    wire new_AGEMA_signal_25357 ;
    wire new_AGEMA_signal_25358 ;
    wire new_AGEMA_signal_25359 ;
    wire new_AGEMA_signal_25360 ;
    wire new_AGEMA_signal_25361 ;
    wire new_AGEMA_signal_25362 ;
    wire new_AGEMA_signal_25363 ;
    wire new_AGEMA_signal_25364 ;
    wire new_AGEMA_signal_25365 ;
    wire new_AGEMA_signal_25366 ;
    wire new_AGEMA_signal_25367 ;
    wire new_AGEMA_signal_25368 ;
    wire new_AGEMA_signal_25369 ;
    wire new_AGEMA_signal_25370 ;
    wire new_AGEMA_signal_25371 ;
    wire new_AGEMA_signal_25372 ;
    wire new_AGEMA_signal_25373 ;
    wire new_AGEMA_signal_25374 ;
    wire new_AGEMA_signal_25375 ;
    wire new_AGEMA_signal_25376 ;
    wire new_AGEMA_signal_25377 ;
    wire new_AGEMA_signal_25378 ;
    wire new_AGEMA_signal_25379 ;
    wire new_AGEMA_signal_25380 ;
    wire new_AGEMA_signal_25381 ;
    wire new_AGEMA_signal_25382 ;
    wire new_AGEMA_signal_25383 ;
    wire new_AGEMA_signal_25384 ;
    wire new_AGEMA_signal_25385 ;
    wire new_AGEMA_signal_25386 ;
    wire new_AGEMA_signal_25387 ;
    wire new_AGEMA_signal_25388 ;
    wire new_AGEMA_signal_25389 ;
    wire new_AGEMA_signal_25390 ;
    wire new_AGEMA_signal_25391 ;
    wire new_AGEMA_signal_25392 ;
    wire new_AGEMA_signal_25393 ;
    wire new_AGEMA_signal_25394 ;
    wire new_AGEMA_signal_25395 ;
    wire new_AGEMA_signal_25396 ;
    wire new_AGEMA_signal_25397 ;
    wire new_AGEMA_signal_25398 ;
    wire new_AGEMA_signal_25399 ;
    wire new_AGEMA_signal_25400 ;
    wire new_AGEMA_signal_25401 ;
    wire new_AGEMA_signal_25402 ;
    wire new_AGEMA_signal_25403 ;
    wire new_AGEMA_signal_25404 ;
    wire new_AGEMA_signal_25405 ;
    wire new_AGEMA_signal_25406 ;
    wire new_AGEMA_signal_25407 ;
    wire new_AGEMA_signal_25408 ;
    wire new_AGEMA_signal_25409 ;
    wire new_AGEMA_signal_25410 ;
    wire new_AGEMA_signal_25411 ;
    wire new_AGEMA_signal_25412 ;
    wire new_AGEMA_signal_25413 ;
    wire new_AGEMA_signal_25414 ;
    wire new_AGEMA_signal_25415 ;
    wire new_AGEMA_signal_25416 ;
    wire new_AGEMA_signal_25417 ;
    wire new_AGEMA_signal_25418 ;
    wire new_AGEMA_signal_25419 ;
    wire new_AGEMA_signal_25420 ;
    wire new_AGEMA_signal_25421 ;
    wire new_AGEMA_signal_25422 ;
    wire new_AGEMA_signal_25423 ;
    wire new_AGEMA_signal_25424 ;
    wire new_AGEMA_signal_25425 ;
    wire new_AGEMA_signal_25426 ;
    wire new_AGEMA_signal_25427 ;
    wire new_AGEMA_signal_25428 ;
    wire new_AGEMA_signal_25429 ;
    wire new_AGEMA_signal_25430 ;
    wire new_AGEMA_signal_25431 ;
    wire new_AGEMA_signal_25432 ;
    wire new_AGEMA_signal_25433 ;
    wire new_AGEMA_signal_25434 ;
    wire new_AGEMA_signal_25435 ;
    wire new_AGEMA_signal_25436 ;
    wire new_AGEMA_signal_25437 ;
    wire new_AGEMA_signal_25438 ;
    wire new_AGEMA_signal_25439 ;
    wire new_AGEMA_signal_25440 ;
    wire new_AGEMA_signal_25441 ;
    wire new_AGEMA_signal_25442 ;
    wire new_AGEMA_signal_25443 ;
    wire new_AGEMA_signal_25444 ;
    wire new_AGEMA_signal_25445 ;
    wire new_AGEMA_signal_25446 ;
    wire new_AGEMA_signal_25447 ;
    wire new_AGEMA_signal_25448 ;
    wire new_AGEMA_signal_25449 ;
    wire new_AGEMA_signal_25450 ;
    wire new_AGEMA_signal_25451 ;
    wire new_AGEMA_signal_25452 ;
    wire new_AGEMA_signal_25453 ;
    wire new_AGEMA_signal_25454 ;
    wire new_AGEMA_signal_25455 ;
    wire new_AGEMA_signal_25456 ;
    wire new_AGEMA_signal_25457 ;
    wire new_AGEMA_signal_25458 ;
    wire new_AGEMA_signal_25459 ;
    wire new_AGEMA_signal_25460 ;
    wire new_AGEMA_signal_25461 ;
    wire new_AGEMA_signal_25462 ;
    wire new_AGEMA_signal_25463 ;
    wire new_AGEMA_signal_25464 ;
    wire new_AGEMA_signal_25465 ;
    wire new_AGEMA_signal_25466 ;
    wire new_AGEMA_signal_25467 ;
    wire new_AGEMA_signal_25468 ;
    wire new_AGEMA_signal_25469 ;
    wire new_AGEMA_signal_25470 ;
    wire new_AGEMA_signal_25471 ;
    wire new_AGEMA_signal_25472 ;
    wire new_AGEMA_signal_25473 ;
    wire new_AGEMA_signal_25474 ;
    wire new_AGEMA_signal_25475 ;
    wire new_AGEMA_signal_25476 ;
    wire new_AGEMA_signal_25477 ;
    wire new_AGEMA_signal_25478 ;
    wire new_AGEMA_signal_25479 ;
    wire new_AGEMA_signal_25480 ;
    wire new_AGEMA_signal_25481 ;
    wire new_AGEMA_signal_25482 ;
    wire new_AGEMA_signal_25483 ;
    wire new_AGEMA_signal_25484 ;
    wire new_AGEMA_signal_25485 ;
    wire new_AGEMA_signal_25486 ;
    wire new_AGEMA_signal_25487 ;
    wire new_AGEMA_signal_25488 ;
    wire new_AGEMA_signal_25489 ;
    wire new_AGEMA_signal_25490 ;
    wire new_AGEMA_signal_25491 ;
    wire new_AGEMA_signal_25492 ;
    wire new_AGEMA_signal_25493 ;
    wire new_AGEMA_signal_25494 ;
    wire new_AGEMA_signal_25495 ;
    wire new_AGEMA_signal_25496 ;
    wire new_AGEMA_signal_25497 ;
    wire new_AGEMA_signal_25498 ;
    wire new_AGEMA_signal_25499 ;
    wire new_AGEMA_signal_25500 ;
    wire new_AGEMA_signal_25501 ;
    wire new_AGEMA_signal_25502 ;
    wire new_AGEMA_signal_25503 ;
    wire new_AGEMA_signal_25504 ;
    wire new_AGEMA_signal_25505 ;
    wire new_AGEMA_signal_25506 ;
    wire new_AGEMA_signal_25507 ;
    wire new_AGEMA_signal_25508 ;
    wire new_AGEMA_signal_25509 ;
    wire new_AGEMA_signal_25510 ;
    wire new_AGEMA_signal_25511 ;
    wire new_AGEMA_signal_25512 ;
    wire new_AGEMA_signal_25513 ;
    wire new_AGEMA_signal_25514 ;
    wire new_AGEMA_signal_25515 ;
    wire new_AGEMA_signal_25516 ;
    wire new_AGEMA_signal_25517 ;
    wire new_AGEMA_signal_25518 ;
    wire new_AGEMA_signal_25519 ;
    wire new_AGEMA_signal_25520 ;
    wire new_AGEMA_signal_25521 ;
    wire new_AGEMA_signal_25522 ;
    wire new_AGEMA_signal_25523 ;
    wire new_AGEMA_signal_25524 ;
    wire new_AGEMA_signal_25525 ;
    wire new_AGEMA_signal_25526 ;
    wire new_AGEMA_signal_25527 ;
    wire new_AGEMA_signal_25528 ;
    wire new_AGEMA_signal_25529 ;
    wire new_AGEMA_signal_25530 ;
    wire new_AGEMA_signal_25531 ;
    wire new_AGEMA_signal_25532 ;
    wire new_AGEMA_signal_25533 ;
    wire new_AGEMA_signal_25534 ;
    wire new_AGEMA_signal_25535 ;
    wire new_AGEMA_signal_25536 ;
    wire new_AGEMA_signal_25537 ;
    wire new_AGEMA_signal_25538 ;
    wire new_AGEMA_signal_25539 ;
    wire new_AGEMA_signal_25540 ;
    wire new_AGEMA_signal_25541 ;
    wire new_AGEMA_signal_25542 ;
    wire new_AGEMA_signal_25543 ;
    wire new_AGEMA_signal_25544 ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U986 ( .a ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U987 ( .a ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, RoundInput[100]}), .b ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, RoundKey[100]}), .c ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U988 ( .a ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundInput[101]}), .b ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, RoundKey[101]}), .c ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U989 ( .a ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[102]}), .b ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, RoundKey[102]}), .c ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U990 ( .a ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, RoundInput[103]}), .b ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, RoundKey[103]}), .c ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U991 ( .a ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundInput[104]}), .b ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, RoundKey[104]}), .c ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U992 ( .a ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[105]}), .b ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, RoundKey[105]}), .c ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U993 ( .a ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, RoundInput[106]}), .b ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, RoundKey[106]}), .c ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U994 ( .a ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundInput[107]}), .b ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, RoundKey[107]}), .c ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U995 ( .a ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[108]}), .b ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, RoundKey[108]}), .c ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U996 ( .a ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, RoundInput[109]}), .b ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, RoundKey[109]}), .c ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U997 ( .a ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundInput[10]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U998 ( .a ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[110]}), .b ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, RoundKey[110]}), .c ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U999 ( .a ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, RoundInput[111]}), .b ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, RoundKey[111]}), .c ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1000 ( .a ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundInput[112]}), .b ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, RoundKey[112]}), .c ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1001 ( .a ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[113]}), .b ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, RoundKey[113]}), .c ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1002 ( .a ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, RoundInput[114]}), .b ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, RoundKey[114]}), .c ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1003 ( .a ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundInput[115]}), .b ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, RoundKey[115]}), .c ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1004 ( .a ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[116]}), .b ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, RoundKey[116]}), .c ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1005 ( .a ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, RoundInput[117]}), .b ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, RoundKey[117]}), .c ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1006 ( .a ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundInput[118]}), .b ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, RoundKey[118]}), .c ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1007 ( .a ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[119]}), .b ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, RoundKey[119]}), .c ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1008 ( .a ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, RoundInput[11]}), .b ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}), .c ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1009 ( .a ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundInput[120]}), .b ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, RoundKey[120]}), .c ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1010 ( .a ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[121]}), .b ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, RoundKey[121]}), .c ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1011 ( .a ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, RoundInput[122]}), .b ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, RoundKey[122]}), .c ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1012 ( .a ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundInput[123]}), .b ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, RoundKey[123]}), .c ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1013 ( .a ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[124]}), .b ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, RoundKey[124]}), .c ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1014 ( .a ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, RoundInput[125]}), .b ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, RoundKey[125]}), .c ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1015 ( .a ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundInput[126]}), .b ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, RoundKey[126]}), .c ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1016 ( .a ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[127]}), .b ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, RoundKey[127]}), .c ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1017 ( .a ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, RoundInput[12]}), .b ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .c ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1018 ( .a ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundInput[13]}), .b ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .c ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1019 ( .a ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[14]}), .b ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .c ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1020 ( .a ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, RoundInput[15]}), .b ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .c ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1021 ( .a ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundInput[16]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1022 ( .a ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[17]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1023 ( .a ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, RoundInput[18]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1024 ( .a ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundInput[19]}), .b ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}), .c ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1025 ( .a ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[1]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1026 ( .a ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, RoundInput[20]}), .b ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .c ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1027 ( .a ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundInput[21]}), .b ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .c ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1028 ( .a ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[22]}), .b ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .c ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1029 ( .a ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, RoundInput[23]}), .b ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .c ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1030 ( .a ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundInput[24]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1031 ( .a ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[25]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1032 ( .a ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, RoundInput[26]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1033 ( .a ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundInput[27]}), .b ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}), .c ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1034 ( .a ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[28]}), .b ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .c ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1035 ( .a ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, RoundInput[29]}), .b ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .c ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1036 ( .a ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundInput[2]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1037 ( .a ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[30]}), .b ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .c ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1038 ( .a ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, RoundInput[31]}), .b ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .c ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1039 ( .a ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundInput[32]}), .b ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, RoundKey[32]}), .c ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1040 ( .a ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[33]}), .b ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, RoundKey[33]}), .c ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1041 ( .a ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, RoundInput[34]}), .b ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, RoundKey[34]}), .c ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1042 ( .a ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundInput[35]}), .b ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, RoundKey[35]}), .c ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1043 ( .a ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[36]}), .b ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, RoundKey[36]}), .c ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1044 ( .a ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, RoundInput[37]}), .b ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, RoundKey[37]}), .c ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1045 ( .a ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundInput[38]}), .b ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, RoundKey[38]}), .c ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1046 ( .a ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[39]}), .b ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, RoundKey[39]}), .c ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1047 ( .a ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, RoundInput[3]}), .b ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}), .c ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1048 ( .a ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundInput[40]}), .b ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, RoundKey[40]}), .c ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1049 ( .a ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[41]}), .b ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, RoundKey[41]}), .c ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1050 ( .a ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, RoundInput[42]}), .b ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, RoundKey[42]}), .c ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1051 ( .a ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundInput[43]}), .b ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, RoundKey[43]}), .c ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1052 ( .a ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[44]}), .b ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, RoundKey[44]}), .c ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1053 ( .a ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, RoundInput[45]}), .b ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, RoundKey[45]}), .c ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1054 ( .a ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundInput[46]}), .b ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, RoundKey[46]}), .c ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1055 ( .a ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[47]}), .b ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, RoundKey[47]}), .c ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1056 ( .a ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, RoundInput[48]}), .b ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, RoundKey[48]}), .c ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1057 ( .a ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundInput[49]}), .b ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, RoundKey[49]}), .c ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1058 ( .a ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[4]}), .b ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .c ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1059 ( .a ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, RoundInput[50]}), .b ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, RoundKey[50]}), .c ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1060 ( .a ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundInput[51]}), .b ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, RoundKey[51]}), .c ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1061 ( .a ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[52]}), .b ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, RoundKey[52]}), .c ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1062 ( .a ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, RoundInput[53]}), .b ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, RoundKey[53]}), .c ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1063 ( .a ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundInput[54]}), .b ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, RoundKey[54]}), .c ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1064 ( .a ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[55]}), .b ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, RoundKey[55]}), .c ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1065 ( .a ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, RoundInput[56]}), .b ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, RoundKey[56]}), .c ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1066 ( .a ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundInput[57]}), .b ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, RoundKey[57]}), .c ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1067 ( .a ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[58]}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, RoundKey[58]}), .c ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1068 ( .a ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, RoundInput[59]}), .b ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, RoundKey[59]}), .c ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1069 ( .a ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundInput[5]}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .c ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1070 ( .a ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[60]}), .b ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, RoundKey[60]}), .c ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1071 ( .a ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, RoundInput[61]}), .b ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, RoundKey[61]}), .c ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1072 ( .a ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundInput[62]}), .b ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, RoundKey[62]}), .c ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1073 ( .a ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[63]}), .b ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, RoundKey[63]}), .c ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1074 ( .a ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, RoundInput[64]}), .b ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, RoundKey[64]}), .c ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1075 ( .a ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundInput[65]}), .b ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, RoundKey[65]}), .c ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1076 ( .a ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[66]}), .b ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, RoundKey[66]}), .c ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1077 ( .a ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, RoundInput[67]}), .b ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, RoundKey[67]}), .c ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1078 ( .a ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundInput[68]}), .b ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, RoundKey[68]}), .c ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1079 ( .a ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[69]}), .b ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, RoundKey[69]}), .c ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1080 ( .a ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, RoundInput[6]}), .b ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .c ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1081 ( .a ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundInput[70]}), .b ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, RoundKey[70]}), .c ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1082 ( .a ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[71]}), .b ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, RoundKey[71]}), .c ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1083 ( .a ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, RoundInput[72]}), .b ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, RoundKey[72]}), .c ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1084 ( .a ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundInput[73]}), .b ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, RoundKey[73]}), .c ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1085 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[74]}), .b ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, RoundKey[74]}), .c ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1086 ( .a ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, RoundInput[75]}), .b ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, RoundKey[75]}), .c ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1087 ( .a ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundInput[76]}), .b ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, RoundKey[76]}), .c ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1088 ( .a ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[77]}), .b ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, RoundKey[77]}), .c ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1089 ( .a ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, RoundInput[78]}), .b ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, RoundKey[78]}), .c ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1090 ( .a ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundInput[79]}), .b ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, RoundKey[79]}), .c ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1091 ( .a ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[7]}), .b ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .c ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1092 ( .a ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, RoundInput[80]}), .b ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, RoundKey[80]}), .c ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1093 ( .a ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundInput[81]}), .b ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, RoundKey[81]}), .c ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1094 ( .a ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[82]}), .b ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, RoundKey[82]}), .c ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1095 ( .a ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, RoundInput[83]}), .b ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, RoundKey[83]}), .c ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1096 ( .a ({new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundInput[84]}), .b ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, RoundKey[84]}), .c ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1097 ( .a ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[85]}), .b ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, RoundKey[85]}), .c ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1098 ( .a ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, RoundInput[86]}), .b ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, RoundKey[86]}), .c ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1099 ( .a ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundInput[87]}), .b ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, RoundKey[87]}), .c ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1100 ( .a ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[88]}), .b ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, RoundKey[88]}), .c ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1101 ( .a ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, RoundInput[89]}), .b ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, RoundKey[89]}), .c ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1102 ( .a ({new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundInput[8]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1103 ( .a ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[90]}), .b ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, RoundKey[90]}), .c ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1104 ( .a ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, RoundInput[91]}), .b ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, RoundKey[91]}), .c ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1105 ( .a ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundInput[92]}), .b ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, RoundKey[92]}), .c ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1106 ( .a ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[93]}), .b ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, RoundKey[93]}), .c ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1107 ( .a ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, RoundInput[94]}), .b ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, RoundKey[94]}), .c ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1108 ( .a ({new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundInput[95]}), .b ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, RoundKey[95]}), .c ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1109 ( .a ({new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[96]}), .b ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, RoundKey[96]}), .c ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1110 ( .a ({new_AGEMA_signal_5294, new_AGEMA_signal_5293, RoundInput[97]}), .b ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, RoundKey[97]}), .c ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1111 ( .a ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundInput[98]}), .b ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, RoundKey[98]}), .c ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1112 ( .a ({new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[99]}), .b ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, RoundKey[99]}), .c ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U1113 ( .a ({new_AGEMA_signal_5312, new_AGEMA_signal_5311, RoundInput[9]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5788, new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5434, new_AGEMA_signal_5433, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5818, new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5476, new_AGEMA_signal_5475, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6232, new_AGEMA_signal_6231, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_6250, new_AGEMA_signal_6249, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5506, new_AGEMA_signal_5505, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5512, new_AGEMA_signal_5511, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_6302, new_AGEMA_signal_6301, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5530, new_AGEMA_signal_5529, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_5536, new_AGEMA_signal_5535, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_6308, new_AGEMA_signal_6307, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_6310, new_AGEMA_signal_6309, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_6328, new_AGEMA_signal_6327, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5547, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_6350, new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_6362, new_AGEMA_signal_6361, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_6380, new_AGEMA_signal_6379, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_6386, new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_6794, new_AGEMA_signal_6793, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_6812, new_AGEMA_signal_6811, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_6830, new_AGEMA_signal_6829, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_6848, new_AGEMA_signal_6847, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_6466, new_AGEMA_signal_6465, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_6484, new_AGEMA_signal_6483, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_6866, new_AGEMA_signal_6865, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_6884, new_AGEMA_signal_6883, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_6902, new_AGEMA_signal_6901, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_6544, new_AGEMA_signal_6543, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .c ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .c ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .b ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .c ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6038, new_AGEMA_signal_6037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}), .c ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .c ({new_AGEMA_signal_5336, new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5336, new_AGEMA_signal_5335, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_6560, new_AGEMA_signal_6559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6050, new_AGEMA_signal_6049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5332, new_AGEMA_signal_5331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .c ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}), .b ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .c ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .b ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .c ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .b ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}), .c ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6068, new_AGEMA_signal_6067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .c ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6074, new_AGEMA_signal_6073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_6578, new_AGEMA_signal_6577, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6076, new_AGEMA_signal_6075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .c ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .c ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .c ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .b ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}), .c ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6094, new_AGEMA_signal_6093, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .c ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_6596, new_AGEMA_signal_6595, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .c ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .c ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .b ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .c ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .b ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}), .c ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .c ({new_AGEMA_signal_5396, new_AGEMA_signal_5395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5396, new_AGEMA_signal_5395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_6614, new_AGEMA_signal_6613, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5781, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6142, new_AGEMA_signal_6141, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_16935, new_AGEMA_signal_16934, new_AGEMA_signal_16933}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_16938, new_AGEMA_signal_16937, new_AGEMA_signal_16936}), .b ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6148, new_AGEMA_signal_6147, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6160, new_AGEMA_signal_6159, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5788, new_AGEMA_signal_5787, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6166, new_AGEMA_signal_6165, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_6646, new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_6646, new_AGEMA_signal_6645, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_6634, new_AGEMA_signal_6633, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_16941, new_AGEMA_signal_16940, new_AGEMA_signal_16939}), .c ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_16944, new_AGEMA_signal_16943, new_AGEMA_signal_16942}), .c ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6178, new_AGEMA_signal_6177, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_16947, new_AGEMA_signal_16946, new_AGEMA_signal_16945}), .b ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6184, new_AGEMA_signal_6183, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5800, new_AGEMA_signal_5799, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_16950, new_AGEMA_signal_16949, new_AGEMA_signal_16948}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_6664, new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_6664, new_AGEMA_signal_6663, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_16953, new_AGEMA_signal_16952, new_AGEMA_signal_16951}), .c ({new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_16956, new_AGEMA_signal_16955, new_AGEMA_signal_16954}), .c ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5818, new_AGEMA_signal_5817, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_16959, new_AGEMA_signal_16958, new_AGEMA_signal_16957}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5824, new_AGEMA_signal_5823, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_16962, new_AGEMA_signal_16961, new_AGEMA_signal_16960}), .b ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6201, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6196, new_AGEMA_signal_6195, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_6682, new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_6682, new_AGEMA_signal_6681, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_16965, new_AGEMA_signal_16964, new_AGEMA_signal_16963}), .c ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6214, new_AGEMA_signal_6213, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_16968, new_AGEMA_signal_16967, new_AGEMA_signal_16966}), .c ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6220, new_AGEMA_signal_6219, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_16971, new_AGEMA_signal_16970, new_AGEMA_signal_16969}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5842, new_AGEMA_signal_5841, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_16974, new_AGEMA_signal_16973, new_AGEMA_signal_16972}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6237, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5836, new_AGEMA_signal_5835, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_6700, new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_6700, new_AGEMA_signal_6699, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_16977, new_AGEMA_signal_16976, new_AGEMA_signal_16975}), .c ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_16980, new_AGEMA_signal_16979, new_AGEMA_signal_16978}), .c ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_6256, new_AGEMA_signal_6255, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_16983, new_AGEMA_signal_16982, new_AGEMA_signal_16981}), .b ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5854, new_AGEMA_signal_5853, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_16986, new_AGEMA_signal_16985, new_AGEMA_signal_16984}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_5860, new_AGEMA_signal_5859, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_6718, new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_6718, new_AGEMA_signal_6717, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_6268, new_AGEMA_signal_6267, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_16989, new_AGEMA_signal_16988, new_AGEMA_signal_16987}), .c ({new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_16992, new_AGEMA_signal_16991, new_AGEMA_signal_16990}), .c ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_16995, new_AGEMA_signal_16994, new_AGEMA_signal_16993}), .b ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_5872, new_AGEMA_signal_5871, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_6286, new_AGEMA_signal_6285, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_16998, new_AGEMA_signal_16997, new_AGEMA_signal_16996}), .b ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6274, new_AGEMA_signal_6273, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_6736, new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_6736, new_AGEMA_signal_6735, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_17001, new_AGEMA_signal_17000, new_AGEMA_signal_16999}), .c ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_6292, new_AGEMA_signal_6291, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_17004, new_AGEMA_signal_17003, new_AGEMA_signal_17002}), .c ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_5878, new_AGEMA_signal_5877, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_6308, new_AGEMA_signal_6307, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_17007, new_AGEMA_signal_17006, new_AGEMA_signal_17005}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_6314, new_AGEMA_signal_6313, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_6314, new_AGEMA_signal_6313, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_5890, new_AGEMA_signal_5889, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_17010, new_AGEMA_signal_17009, new_AGEMA_signal_17008}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_6304, new_AGEMA_signal_6303, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_6322, new_AGEMA_signal_6321, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_6754, new_AGEMA_signal_6753, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_6754, new_AGEMA_signal_6753, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_6320, new_AGEMA_signal_6319, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_17013, new_AGEMA_signal_17012, new_AGEMA_signal_17011}), .c ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_17016, new_AGEMA_signal_17015, new_AGEMA_signal_17014}), .c ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_17019, new_AGEMA_signal_17018, new_AGEMA_signal_17017}), .b ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_6340, new_AGEMA_signal_6339, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_6338, new_AGEMA_signal_6337, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_5896, new_AGEMA_signal_5895, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_6344, new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_17022, new_AGEMA_signal_17021, new_AGEMA_signal_17020}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_6332, new_AGEMA_signal_6331, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6325, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_6772, new_AGEMA_signal_6771, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_6772, new_AGEMA_signal_6771, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_6346, new_AGEMA_signal_6345, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_17025, new_AGEMA_signal_17024, new_AGEMA_signal_17023}), .c ({new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_6344, new_AGEMA_signal_6343, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_17028, new_AGEMA_signal_17027, new_AGEMA_signal_17026}), .c ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_6350, new_AGEMA_signal_6349, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_17031, new_AGEMA_signal_17030, new_AGEMA_signal_17029}), .b ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_6364, new_AGEMA_signal_6363, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_6782, new_AGEMA_signal_6781, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_17034, new_AGEMA_signal_17033, new_AGEMA_signal_17032}), .b ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6357, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_6356, new_AGEMA_signal_6355, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_6368, new_AGEMA_signal_6367, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_6374, new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_6374, new_AGEMA_signal_6373, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_6790, new_AGEMA_signal_6789, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_6790, new_AGEMA_signal_6789, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_6782, new_AGEMA_signal_6781, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_17037, new_AGEMA_signal_17036, new_AGEMA_signal_17035}), .c ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_6788, new_AGEMA_signal_6787, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_17040, new_AGEMA_signal_17039, new_AGEMA_signal_17038}), .c ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5925, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_6386, new_AGEMA_signal_6385, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_6376, new_AGEMA_signal_6375, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_6796, new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_17043, new_AGEMA_signal_17042, new_AGEMA_signal_17041}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_6392, new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_6392, new_AGEMA_signal_6391, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_6800, new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_17046, new_AGEMA_signal_17045, new_AGEMA_signal_17044}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_6382, new_AGEMA_signal_6381, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6393, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_5932, new_AGEMA_signal_5931, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_6400, new_AGEMA_signal_6399, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_6808, new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_6808, new_AGEMA_signal_6807, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_6796, new_AGEMA_signal_6795, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_6800, new_AGEMA_signal_6799, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_17049, new_AGEMA_signal_17048, new_AGEMA_signal_17047}), .c ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6805, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_17052, new_AGEMA_signal_17051, new_AGEMA_signal_17050}), .c ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_7568, new_AGEMA_signal_7567, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_6412, new_AGEMA_signal_6411, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_6814, new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_17055, new_AGEMA_signal_17054, new_AGEMA_signal_17053}), .b ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_6418, new_AGEMA_signal_6417, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_6818, new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_5950, new_AGEMA_signal_5949, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_5944, new_AGEMA_signal_5943, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_17058, new_AGEMA_signal_17057, new_AGEMA_signal_17056}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_6826, new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_6826, new_AGEMA_signal_6825, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_6814, new_AGEMA_signal_6813, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_6818, new_AGEMA_signal_6817, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_17061, new_AGEMA_signal_17060, new_AGEMA_signal_17059}), .c ({new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_6824, new_AGEMA_signal_6823, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_17064, new_AGEMA_signal_17063, new_AGEMA_signal_17062}), .c ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_5962, new_AGEMA_signal_5961, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_6832, new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_17067, new_AGEMA_signal_17066, new_AGEMA_signal_17065}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_5968, new_AGEMA_signal_5967, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_6836, new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_17070, new_AGEMA_signal_17069, new_AGEMA_signal_17068}), .b ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_6436, new_AGEMA_signal_6435, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6429, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_6844, new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_6844, new_AGEMA_signal_6843, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_6832, new_AGEMA_signal_6831, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_6836, new_AGEMA_signal_6835, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_17073, new_AGEMA_signal_17072, new_AGEMA_signal_17071}), .c ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_6448, new_AGEMA_signal_6447, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_6842, new_AGEMA_signal_6841, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_17076, new_AGEMA_signal_17075, new_AGEMA_signal_17074}), .c ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_6454, new_AGEMA_signal_6453, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_6850, new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_17079, new_AGEMA_signal_17078, new_AGEMA_signal_17077}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_6854, new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_5986, new_AGEMA_signal_5985, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_17082, new_AGEMA_signal_17081, new_AGEMA_signal_17080}), .b ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_6472, new_AGEMA_signal_6471, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_5980, new_AGEMA_signal_5979, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_6862, new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_6862, new_AGEMA_signal_6861, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_6850, new_AGEMA_signal_6849, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_6854, new_AGEMA_signal_6853, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_17085, new_AGEMA_signal_17084, new_AGEMA_signal_17083}), .c ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_6860, new_AGEMA_signal_6859, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_17088, new_AGEMA_signal_17087, new_AGEMA_signal_17086}), .c ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_7598, new_AGEMA_signal_7597, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_6490, new_AGEMA_signal_6489, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_6868, new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_17091, new_AGEMA_signal_17090, new_AGEMA_signal_17089}), .b ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_6872, new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5997, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_17094, new_AGEMA_signal_17093, new_AGEMA_signal_17092}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_6004, new_AGEMA_signal_6003, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_6880, new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_6880, new_AGEMA_signal_6879, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_6502, new_AGEMA_signal_6501, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_6868, new_AGEMA_signal_6867, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_6872, new_AGEMA_signal_6871, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_17097, new_AGEMA_signal_17096, new_AGEMA_signal_17095}), .c ({new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_6878, new_AGEMA_signal_6877, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_17100, new_AGEMA_signal_17099, new_AGEMA_signal_17098}), .c ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_17103, new_AGEMA_signal_17102, new_AGEMA_signal_17101}), .b ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_6016, new_AGEMA_signal_6015, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_6520, new_AGEMA_signal_6519, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_6890, new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_17106, new_AGEMA_signal_17105, new_AGEMA_signal_17104}), .b ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6508, new_AGEMA_signal_6507, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_6890, new_AGEMA_signal_6889, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_17109, new_AGEMA_signal_17108, new_AGEMA_signal_17107}), .c ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_6526, new_AGEMA_signal_6525, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_6896, new_AGEMA_signal_6895, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_17112, new_AGEMA_signal_17111, new_AGEMA_signal_17110}), .c ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_6022, new_AGEMA_signal_6021, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_17115, new_AGEMA_signal_17114, new_AGEMA_signal_17113}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_6908, new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_6034, new_AGEMA_signal_6033, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_17118, new_AGEMA_signal_17117, new_AGEMA_signal_17116}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6537, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_6556, new_AGEMA_signal_6555, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_6556, new_AGEMA_signal_6555, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_6908, new_AGEMA_signal_6907, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_17121, new_AGEMA_signal_17120, new_AGEMA_signal_17119}), .c ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_6914, new_AGEMA_signal_6913, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_17124, new_AGEMA_signal_17123, new_AGEMA_signal_17122}), .c ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_7628, new_AGEMA_signal_7627, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6038, new_AGEMA_signal_6037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_6562, new_AGEMA_signal_6561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_17127, new_AGEMA_signal_17126, new_AGEMA_signal_17125}), .b ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6052, new_AGEMA_signal_6051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_6566, new_AGEMA_signal_6565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_17130, new_AGEMA_signal_17129, new_AGEMA_signal_17128}), .b ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6044, new_AGEMA_signal_6043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6056, new_AGEMA_signal_6055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_6062, new_AGEMA_signal_6061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6062, new_AGEMA_signal_6061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5320, new_AGEMA_signal_5319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6040, new_AGEMA_signal_6039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_6574, new_AGEMA_signal_6573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_6562, new_AGEMA_signal_6561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_6566, new_AGEMA_signal_6565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_17133, new_AGEMA_signal_17132, new_AGEMA_signal_17131}), .c ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6058, new_AGEMA_signal_6057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_6572, new_AGEMA_signal_6571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_17136, new_AGEMA_signal_17135, new_AGEMA_signal_17134}), .c ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6074, new_AGEMA_signal_6073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_17139, new_AGEMA_signal_17138, new_AGEMA_signal_17137}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_6080, new_AGEMA_signal_6079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6080, new_AGEMA_signal_6079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5342, new_AGEMA_signal_5341, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_17142, new_AGEMA_signal_17141, new_AGEMA_signal_17140}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6070, new_AGEMA_signal_6069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6088, new_AGEMA_signal_6087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_6592, new_AGEMA_signal_6591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6086, new_AGEMA_signal_6085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_6580, new_AGEMA_signal_6579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_17145, new_AGEMA_signal_17144, new_AGEMA_signal_17143}), .c ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_17148, new_AGEMA_signal_17147, new_AGEMA_signal_17146}), .c ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_7448, new_AGEMA_signal_7447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_17151, new_AGEMA_signal_17150, new_AGEMA_signal_17149}), .b ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6106, new_AGEMA_signal_6105, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_17154, new_AGEMA_signal_17153, new_AGEMA_signal_17152}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_6938, new_AGEMA_signal_6937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5360, new_AGEMA_signal_5359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_6610, new_AGEMA_signal_6609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6112, new_AGEMA_signal_6111, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_6598, new_AGEMA_signal_6597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_17157, new_AGEMA_signal_17156, new_AGEMA_signal_17155}), .c ({new_AGEMA_signal_6944, new_AGEMA_signal_6943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_6938, new_AGEMA_signal_6937, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_6944, new_AGEMA_signal_6943, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_17160, new_AGEMA_signal_17159, new_AGEMA_signal_17158}), .c ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_7298, new_AGEMA_signal_7297, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_17163, new_AGEMA_signal_17162, new_AGEMA_signal_17161}), .b ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6130, new_AGEMA_signal_6129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_17166, new_AGEMA_signal_17165, new_AGEMA_signal_17164}), .b ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6124, new_AGEMA_signal_6123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5384, new_AGEMA_signal_5383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_6628, new_AGEMA_signal_6627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_6616, new_AGEMA_signal_6615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_17169, new_AGEMA_signal_17168, new_AGEMA_signal_17167}), .c ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_6956, new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_6950, new_AGEMA_signal_6949, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_6956, new_AGEMA_signal_6955, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_17172, new_AGEMA_signal_17171, new_AGEMA_signal_17170}), .c ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_16933) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_6145), .Q (new_AGEMA_signal_16934) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_16935) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_16936) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_16937) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_16938) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_16939) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_6629), .Q (new_AGEMA_signal_16940) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_16941) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_16942) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_16943) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_16944) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_16945) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_16946) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_16947) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_16948) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_16949) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_16950) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_16951) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_16952) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_16953) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_16954) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_16955) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_6650), .Q (new_AGEMA_signal_16956) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_16957) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_6197), .Q (new_AGEMA_signal_16958) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_16959) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_16960) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_6205), .Q (new_AGEMA_signal_16961) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_16962) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_16963) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_6665), .Q (new_AGEMA_signal_16964) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_6666), .Q (new_AGEMA_signal_16965) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_16966) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_16967) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_16968) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_16969) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_16970) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_16971) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_16972) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_16973) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_16974) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_16975) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_16976) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_16977) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_16978) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_16979) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_6686), .Q (new_AGEMA_signal_16980) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T14), .Q (new_AGEMA_signal_16981) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_16982) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_16983) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T26), .Q (new_AGEMA_signal_16984) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_6257), .Q (new_AGEMA_signal_16985) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_16986) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T24), .Q (new_AGEMA_signal_16987) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_6701), .Q (new_AGEMA_signal_16988) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_16989) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T25), .Q (new_AGEMA_signal_16990) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_16991) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_16992) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T14), .Q (new_AGEMA_signal_16993) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_16994) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_16995) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T26), .Q (new_AGEMA_signal_16996) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_16997) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_16998) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T24), .Q (new_AGEMA_signal_16999) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_17000) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_17001) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T25), .Q (new_AGEMA_signal_17002) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_17003) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_6722), .Q (new_AGEMA_signal_17004) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T14), .Q (new_AGEMA_signal_17005) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_6301), .Q (new_AGEMA_signal_17006) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_17007) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T26), .Q (new_AGEMA_signal_17008) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_17009) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_17010) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T24), .Q (new_AGEMA_signal_17011) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_6737), .Q (new_AGEMA_signal_17012) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_6738), .Q (new_AGEMA_signal_17013) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T25), .Q (new_AGEMA_signal_17014) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_17015) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_17016) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T14), .Q (new_AGEMA_signal_17017) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_17018) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_17019) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T26), .Q (new_AGEMA_signal_17020) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_17021) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_17022) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T24), .Q (new_AGEMA_signal_17023) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_17024) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_17025) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T25), .Q (new_AGEMA_signal_17026) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_17027) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_6758), .Q (new_AGEMA_signal_17028) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T14), .Q (new_AGEMA_signal_17029) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_6353), .Q (new_AGEMA_signal_17030) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_17031) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T26), .Q (new_AGEMA_signal_17032) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_6361), .Q (new_AGEMA_signal_17033) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_17034) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T24), .Q (new_AGEMA_signal_17035) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_6773), .Q (new_AGEMA_signal_17036) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_17037) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T25), .Q (new_AGEMA_signal_17038) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_17039) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_17040) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T14), .Q (new_AGEMA_signal_17041) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_17042) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_17043) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T26), .Q (new_AGEMA_signal_17044) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_17045) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_17046) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T24), .Q (new_AGEMA_signal_17047) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_17048) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_17049) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T25), .Q (new_AGEMA_signal_17050) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_17051) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_6794), .Q (new_AGEMA_signal_17052) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T14), .Q (new_AGEMA_signal_17053) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_17054) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_17055) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T26), .Q (new_AGEMA_signal_17056) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_6413), .Q (new_AGEMA_signal_17057) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_17058) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T24), .Q (new_AGEMA_signal_17059) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_6809), .Q (new_AGEMA_signal_17060) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (new_AGEMA_signal_6810), .Q (new_AGEMA_signal_17061) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T25), .Q (new_AGEMA_signal_17062) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_17063) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_17064) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T14), .Q (new_AGEMA_signal_17065) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_17066) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_17067) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T26), .Q (new_AGEMA_signal_17068) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_17069) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_17070) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T24), .Q (new_AGEMA_signal_17071) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_17072) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_17073) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T25), .Q (new_AGEMA_signal_17074) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_6829), .Q (new_AGEMA_signal_17075) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_17076) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T14), .Q (new_AGEMA_signal_17077) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_17078) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_17079) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T26), .Q (new_AGEMA_signal_17080) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_17081) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_17082) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T24), .Q (new_AGEMA_signal_17083) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_6845), .Q (new_AGEMA_signal_17084) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (new_AGEMA_signal_6846), .Q (new_AGEMA_signal_17085) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T25), .Q (new_AGEMA_signal_17086) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_17087) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_17088) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T14), .Q (new_AGEMA_signal_17089) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_17090) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_17091) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T26), .Q (new_AGEMA_signal_17092) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_17093) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_17094) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T24), .Q (new_AGEMA_signal_17095) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_17096) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_17097) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T25), .Q (new_AGEMA_signal_17098) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_6865), .Q (new_AGEMA_signal_17099) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_6866), .Q (new_AGEMA_signal_17100) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T14), .Q (new_AGEMA_signal_17101) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_17102) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_17103) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T26), .Q (new_AGEMA_signal_17104) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (new_AGEMA_signal_6517), .Q (new_AGEMA_signal_17105) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_17106) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T24), .Q (new_AGEMA_signal_17107) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_6881), .Q (new_AGEMA_signal_17108) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (new_AGEMA_signal_6882), .Q (new_AGEMA_signal_17109) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T25), .Q (new_AGEMA_signal_17110) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_17111) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_17112) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T14), .Q (new_AGEMA_signal_17113) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_17114) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_17115) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T26), .Q (new_AGEMA_signal_17116) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_17117) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_17118) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T24), .Q (new_AGEMA_signal_17119) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_17120) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_17121) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T25), .Q (new_AGEMA_signal_17122) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_6901), .Q (new_AGEMA_signal_17123) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_17124) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_17125) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_17126) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_17127) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_17128) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_6049), .Q (new_AGEMA_signal_17129) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_17130) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_17131) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_6557), .Q (new_AGEMA_signal_17132) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_17133) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_17134) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_17135) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_17136) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_17137) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_17138) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_17139) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_17140) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_17141) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_17142) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_17143) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_17144) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_17145) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_17146) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_6577), .Q (new_AGEMA_signal_17147) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_17148) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_17149) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_17150) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_17151) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_17152) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (new_AGEMA_signal_6101), .Q (new_AGEMA_signal_17153) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_17154) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_17155) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_6593), .Q (new_AGEMA_signal_17156) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_17157) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_17158) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_17159) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_17160) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_17161) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_17162) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_17163) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_17164) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_17165) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_17166) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_17167) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_17168) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_17169) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_17170) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_6613), .Q (new_AGEMA_signal_17171) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_17172) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C (clk), .D (n321), .Q (new_AGEMA_signal_17653) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C (clk), .D (n315), .Q (new_AGEMA_signal_17657) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C (clk), .D (n316), .Q (new_AGEMA_signal_17661) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C (clk), .D (n317), .Q (new_AGEMA_signal_17665) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C (clk), .D (n318), .Q (new_AGEMA_signal_17669) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C (clk), .D (n319), .Q (new_AGEMA_signal_17673) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C (clk), .D (n320), .Q (new_AGEMA_signal_17677) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_17681) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_17685) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_17689) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C (clk), .D (plaintext_s2[0]), .Q (new_AGEMA_signal_17693) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_17697) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_17701) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C (clk), .D (plaintext_s2[1]), .Q (new_AGEMA_signal_17705) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_17709) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_17713) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C (clk), .D (plaintext_s2[2]), .Q (new_AGEMA_signal_17717) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_17721) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_17725) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C (clk), .D (plaintext_s2[3]), .Q (new_AGEMA_signal_17729) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_17733) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_17737) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C (clk), .D (plaintext_s2[4]), .Q (new_AGEMA_signal_17741) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_17745) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_17749) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C (clk), .D (plaintext_s2[5]), .Q (new_AGEMA_signal_17753) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_17757) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_17761) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C (clk), .D (plaintext_s2[6]), .Q (new_AGEMA_signal_17765) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_17769) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_17773) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C (clk), .D (plaintext_s2[7]), .Q (new_AGEMA_signal_17777) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_17781) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_17785) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C (clk), .D (plaintext_s2[8]), .Q (new_AGEMA_signal_17789) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_17793) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_17797) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C (clk), .D (plaintext_s2[9]), .Q (new_AGEMA_signal_17801) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_17805) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_17809) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C (clk), .D (plaintext_s2[10]), .Q (new_AGEMA_signal_17813) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_17817) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_17821) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C (clk), .D (plaintext_s2[11]), .Q (new_AGEMA_signal_17825) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_17829) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_17833) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C (clk), .D (plaintext_s2[12]), .Q (new_AGEMA_signal_17837) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_17841) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_17845) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C (clk), .D (plaintext_s2[13]), .Q (new_AGEMA_signal_17849) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_17853) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_17857) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C (clk), .D (plaintext_s2[14]), .Q (new_AGEMA_signal_17861) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_17865) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_17869) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C (clk), .D (plaintext_s2[15]), .Q (new_AGEMA_signal_17873) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_17877) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_17881) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C (clk), .D (plaintext_s2[16]), .Q (new_AGEMA_signal_17885) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_17889) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_17893) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C (clk), .D (plaintext_s2[17]), .Q (new_AGEMA_signal_17897) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_17901) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_17905) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C (clk), .D (plaintext_s2[18]), .Q (new_AGEMA_signal_17909) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_17913) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_17917) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C (clk), .D (plaintext_s2[19]), .Q (new_AGEMA_signal_17921) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_17925) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_17929) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C (clk), .D (plaintext_s2[20]), .Q (new_AGEMA_signal_17933) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_17937) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_17941) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C (clk), .D (plaintext_s2[21]), .Q (new_AGEMA_signal_17945) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_17949) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_17953) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C (clk), .D (plaintext_s2[22]), .Q (new_AGEMA_signal_17957) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_17961) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_17965) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C (clk), .D (plaintext_s2[23]), .Q (new_AGEMA_signal_17969) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_17973) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_17977) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C (clk), .D (plaintext_s2[24]), .Q (new_AGEMA_signal_17981) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_17985) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_17989) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C (clk), .D (plaintext_s2[25]), .Q (new_AGEMA_signal_17993) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_17997) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_18001) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C (clk), .D (plaintext_s2[26]), .Q (new_AGEMA_signal_18005) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_18009) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_18013) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C (clk), .D (plaintext_s2[27]), .Q (new_AGEMA_signal_18017) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_18021) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_18025) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C (clk), .D (plaintext_s2[28]), .Q (new_AGEMA_signal_18029) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_18033) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_18037) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C (clk), .D (plaintext_s2[29]), .Q (new_AGEMA_signal_18041) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_18045) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_18049) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C (clk), .D (plaintext_s2[30]), .Q (new_AGEMA_signal_18053) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_18057) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_18061) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C (clk), .D (plaintext_s2[31]), .Q (new_AGEMA_signal_18065) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_18069) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_18073) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C (clk), .D (plaintext_s2[32]), .Q (new_AGEMA_signal_18077) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_18081) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_18085) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C (clk), .D (plaintext_s2[33]), .Q (new_AGEMA_signal_18089) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_18093) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_18097) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C (clk), .D (plaintext_s2[34]), .Q (new_AGEMA_signal_18101) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_18105) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_18109) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C (clk), .D (plaintext_s2[35]), .Q (new_AGEMA_signal_18113) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_18117) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_18121) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C (clk), .D (plaintext_s2[36]), .Q (new_AGEMA_signal_18125) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_18129) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_18133) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C (clk), .D (plaintext_s2[37]), .Q (new_AGEMA_signal_18137) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_18141) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_18145) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C (clk), .D (plaintext_s2[38]), .Q (new_AGEMA_signal_18149) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_18153) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_18157) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C (clk), .D (plaintext_s2[39]), .Q (new_AGEMA_signal_18161) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_18165) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_18169) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C (clk), .D (plaintext_s2[40]), .Q (new_AGEMA_signal_18173) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_18177) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_18181) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C (clk), .D (plaintext_s2[41]), .Q (new_AGEMA_signal_18185) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_18189) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_18193) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C (clk), .D (plaintext_s2[42]), .Q (new_AGEMA_signal_18197) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_18201) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_18205) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C (clk), .D (plaintext_s2[43]), .Q (new_AGEMA_signal_18209) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_18213) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_18217) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C (clk), .D (plaintext_s2[44]), .Q (new_AGEMA_signal_18221) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_18225) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_18229) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C (clk), .D (plaintext_s2[45]), .Q (new_AGEMA_signal_18233) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_18237) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_18241) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C (clk), .D (plaintext_s2[46]), .Q (new_AGEMA_signal_18245) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_18249) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_18253) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C (clk), .D (plaintext_s2[47]), .Q (new_AGEMA_signal_18257) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_18261) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_18265) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C (clk), .D (plaintext_s2[48]), .Q (new_AGEMA_signal_18269) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_18273) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_18277) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C (clk), .D (plaintext_s2[49]), .Q (new_AGEMA_signal_18281) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_18285) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_18289) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C (clk), .D (plaintext_s2[50]), .Q (new_AGEMA_signal_18293) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_18297) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_18301) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C (clk), .D (plaintext_s2[51]), .Q (new_AGEMA_signal_18305) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_18309) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_18313) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C (clk), .D (plaintext_s2[52]), .Q (new_AGEMA_signal_18317) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_18321) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_18325) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C (clk), .D (plaintext_s2[53]), .Q (new_AGEMA_signal_18329) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_18333) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_18337) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C (clk), .D (plaintext_s2[54]), .Q (new_AGEMA_signal_18341) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_18345) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_18349) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C (clk), .D (plaintext_s2[55]), .Q (new_AGEMA_signal_18353) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_18357) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_18361) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C (clk), .D (plaintext_s2[56]), .Q (new_AGEMA_signal_18365) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_18369) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_18373) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C (clk), .D (plaintext_s2[57]), .Q (new_AGEMA_signal_18377) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_18381) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_18385) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C (clk), .D (plaintext_s2[58]), .Q (new_AGEMA_signal_18389) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_18393) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_18397) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C (clk), .D (plaintext_s2[59]), .Q (new_AGEMA_signal_18401) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_18405) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_18409) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C (clk), .D (plaintext_s2[60]), .Q (new_AGEMA_signal_18413) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_18417) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_18421) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C (clk), .D (plaintext_s2[61]), .Q (new_AGEMA_signal_18425) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_18429) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_18433) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C (clk), .D (plaintext_s2[62]), .Q (new_AGEMA_signal_18437) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_18441) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_18445) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C (clk), .D (plaintext_s2[63]), .Q (new_AGEMA_signal_18449) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C (clk), .D (plaintext_s0[64]), .Q (new_AGEMA_signal_18453) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C (clk), .D (plaintext_s1[64]), .Q (new_AGEMA_signal_18457) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C (clk), .D (plaintext_s2[64]), .Q (new_AGEMA_signal_18461) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C (clk), .D (plaintext_s0[65]), .Q (new_AGEMA_signal_18465) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C (clk), .D (plaintext_s1[65]), .Q (new_AGEMA_signal_18469) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C (clk), .D (plaintext_s2[65]), .Q (new_AGEMA_signal_18473) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C (clk), .D (plaintext_s0[66]), .Q (new_AGEMA_signal_18477) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C (clk), .D (plaintext_s1[66]), .Q (new_AGEMA_signal_18481) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C (clk), .D (plaintext_s2[66]), .Q (new_AGEMA_signal_18485) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C (clk), .D (plaintext_s0[67]), .Q (new_AGEMA_signal_18489) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C (clk), .D (plaintext_s1[67]), .Q (new_AGEMA_signal_18493) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C (clk), .D (plaintext_s2[67]), .Q (new_AGEMA_signal_18497) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C (clk), .D (plaintext_s0[68]), .Q (new_AGEMA_signal_18501) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C (clk), .D (plaintext_s1[68]), .Q (new_AGEMA_signal_18505) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C (clk), .D (plaintext_s2[68]), .Q (new_AGEMA_signal_18509) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C (clk), .D (plaintext_s0[69]), .Q (new_AGEMA_signal_18513) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C (clk), .D (plaintext_s1[69]), .Q (new_AGEMA_signal_18517) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C (clk), .D (plaintext_s2[69]), .Q (new_AGEMA_signal_18521) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C (clk), .D (plaintext_s0[70]), .Q (new_AGEMA_signal_18525) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C (clk), .D (plaintext_s1[70]), .Q (new_AGEMA_signal_18529) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C (clk), .D (plaintext_s2[70]), .Q (new_AGEMA_signal_18533) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C (clk), .D (plaintext_s0[71]), .Q (new_AGEMA_signal_18537) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C (clk), .D (plaintext_s1[71]), .Q (new_AGEMA_signal_18541) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C (clk), .D (plaintext_s2[71]), .Q (new_AGEMA_signal_18545) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C (clk), .D (plaintext_s0[72]), .Q (new_AGEMA_signal_18549) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C (clk), .D (plaintext_s1[72]), .Q (new_AGEMA_signal_18553) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C (clk), .D (plaintext_s2[72]), .Q (new_AGEMA_signal_18557) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C (clk), .D (plaintext_s0[73]), .Q (new_AGEMA_signal_18561) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C (clk), .D (plaintext_s1[73]), .Q (new_AGEMA_signal_18565) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C (clk), .D (plaintext_s2[73]), .Q (new_AGEMA_signal_18569) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C (clk), .D (plaintext_s0[74]), .Q (new_AGEMA_signal_18573) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C (clk), .D (plaintext_s1[74]), .Q (new_AGEMA_signal_18577) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C (clk), .D (plaintext_s2[74]), .Q (new_AGEMA_signal_18581) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C (clk), .D (plaintext_s0[75]), .Q (new_AGEMA_signal_18585) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C (clk), .D (plaintext_s1[75]), .Q (new_AGEMA_signal_18589) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C (clk), .D (plaintext_s2[75]), .Q (new_AGEMA_signal_18593) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C (clk), .D (plaintext_s0[76]), .Q (new_AGEMA_signal_18597) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C (clk), .D (plaintext_s1[76]), .Q (new_AGEMA_signal_18601) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C (clk), .D (plaintext_s2[76]), .Q (new_AGEMA_signal_18605) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C (clk), .D (plaintext_s0[77]), .Q (new_AGEMA_signal_18609) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C (clk), .D (plaintext_s1[77]), .Q (new_AGEMA_signal_18613) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C (clk), .D (plaintext_s2[77]), .Q (new_AGEMA_signal_18617) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C (clk), .D (plaintext_s0[78]), .Q (new_AGEMA_signal_18621) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C (clk), .D (plaintext_s1[78]), .Q (new_AGEMA_signal_18625) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C (clk), .D (plaintext_s2[78]), .Q (new_AGEMA_signal_18629) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C (clk), .D (plaintext_s0[79]), .Q (new_AGEMA_signal_18633) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C (clk), .D (plaintext_s1[79]), .Q (new_AGEMA_signal_18637) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C (clk), .D (plaintext_s2[79]), .Q (new_AGEMA_signal_18641) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C (clk), .D (plaintext_s0[80]), .Q (new_AGEMA_signal_18645) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C (clk), .D (plaintext_s1[80]), .Q (new_AGEMA_signal_18649) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C (clk), .D (plaintext_s2[80]), .Q (new_AGEMA_signal_18653) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C (clk), .D (plaintext_s0[81]), .Q (new_AGEMA_signal_18657) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C (clk), .D (plaintext_s1[81]), .Q (new_AGEMA_signal_18661) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C (clk), .D (plaintext_s2[81]), .Q (new_AGEMA_signal_18665) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C (clk), .D (plaintext_s0[82]), .Q (new_AGEMA_signal_18669) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C (clk), .D (plaintext_s1[82]), .Q (new_AGEMA_signal_18673) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C (clk), .D (plaintext_s2[82]), .Q (new_AGEMA_signal_18677) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C (clk), .D (plaintext_s0[83]), .Q (new_AGEMA_signal_18681) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C (clk), .D (plaintext_s1[83]), .Q (new_AGEMA_signal_18685) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C (clk), .D (plaintext_s2[83]), .Q (new_AGEMA_signal_18689) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C (clk), .D (plaintext_s0[84]), .Q (new_AGEMA_signal_18693) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C (clk), .D (plaintext_s1[84]), .Q (new_AGEMA_signal_18697) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C (clk), .D (plaintext_s2[84]), .Q (new_AGEMA_signal_18701) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C (clk), .D (plaintext_s0[85]), .Q (new_AGEMA_signal_18705) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C (clk), .D (plaintext_s1[85]), .Q (new_AGEMA_signal_18709) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C (clk), .D (plaintext_s2[85]), .Q (new_AGEMA_signal_18713) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C (clk), .D (plaintext_s0[86]), .Q (new_AGEMA_signal_18717) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C (clk), .D (plaintext_s1[86]), .Q (new_AGEMA_signal_18721) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C (clk), .D (plaintext_s2[86]), .Q (new_AGEMA_signal_18725) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C (clk), .D (plaintext_s0[87]), .Q (new_AGEMA_signal_18729) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C (clk), .D (plaintext_s1[87]), .Q (new_AGEMA_signal_18733) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C (clk), .D (plaintext_s2[87]), .Q (new_AGEMA_signal_18737) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C (clk), .D (plaintext_s0[88]), .Q (new_AGEMA_signal_18741) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C (clk), .D (plaintext_s1[88]), .Q (new_AGEMA_signal_18745) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C (clk), .D (plaintext_s2[88]), .Q (new_AGEMA_signal_18749) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C (clk), .D (plaintext_s0[89]), .Q (new_AGEMA_signal_18753) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C (clk), .D (plaintext_s1[89]), .Q (new_AGEMA_signal_18757) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C (clk), .D (plaintext_s2[89]), .Q (new_AGEMA_signal_18761) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C (clk), .D (plaintext_s0[90]), .Q (new_AGEMA_signal_18765) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C (clk), .D (plaintext_s1[90]), .Q (new_AGEMA_signal_18769) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C (clk), .D (plaintext_s2[90]), .Q (new_AGEMA_signal_18773) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C (clk), .D (plaintext_s0[91]), .Q (new_AGEMA_signal_18777) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C (clk), .D (plaintext_s1[91]), .Q (new_AGEMA_signal_18781) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C (clk), .D (plaintext_s2[91]), .Q (new_AGEMA_signal_18785) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C (clk), .D (plaintext_s0[92]), .Q (new_AGEMA_signal_18789) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C (clk), .D (plaintext_s1[92]), .Q (new_AGEMA_signal_18793) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C (clk), .D (plaintext_s2[92]), .Q (new_AGEMA_signal_18797) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C (clk), .D (plaintext_s0[93]), .Q (new_AGEMA_signal_18801) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C (clk), .D (plaintext_s1[93]), .Q (new_AGEMA_signal_18805) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C (clk), .D (plaintext_s2[93]), .Q (new_AGEMA_signal_18809) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C (clk), .D (plaintext_s0[94]), .Q (new_AGEMA_signal_18813) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C (clk), .D (plaintext_s1[94]), .Q (new_AGEMA_signal_18817) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C (clk), .D (plaintext_s2[94]), .Q (new_AGEMA_signal_18821) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C (clk), .D (plaintext_s0[95]), .Q (new_AGEMA_signal_18825) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C (clk), .D (plaintext_s1[95]), .Q (new_AGEMA_signal_18829) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C (clk), .D (plaintext_s2[95]), .Q (new_AGEMA_signal_18833) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C (clk), .D (plaintext_s0[96]), .Q (new_AGEMA_signal_18837) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C (clk), .D (plaintext_s1[96]), .Q (new_AGEMA_signal_18841) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C (clk), .D (plaintext_s2[96]), .Q (new_AGEMA_signal_18845) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C (clk), .D (plaintext_s0[97]), .Q (new_AGEMA_signal_18849) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C (clk), .D (plaintext_s1[97]), .Q (new_AGEMA_signal_18853) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C (clk), .D (plaintext_s2[97]), .Q (new_AGEMA_signal_18857) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C (clk), .D (plaintext_s0[98]), .Q (new_AGEMA_signal_18861) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C (clk), .D (plaintext_s1[98]), .Q (new_AGEMA_signal_18865) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C (clk), .D (plaintext_s2[98]), .Q (new_AGEMA_signal_18869) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C (clk), .D (plaintext_s0[99]), .Q (new_AGEMA_signal_18873) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C (clk), .D (plaintext_s1[99]), .Q (new_AGEMA_signal_18877) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C (clk), .D (plaintext_s2[99]), .Q (new_AGEMA_signal_18881) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C (clk), .D (plaintext_s0[100]), .Q (new_AGEMA_signal_18885) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C (clk), .D (plaintext_s1[100]), .Q (new_AGEMA_signal_18889) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C (clk), .D (plaintext_s2[100]), .Q (new_AGEMA_signal_18893) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C (clk), .D (plaintext_s0[101]), .Q (new_AGEMA_signal_18897) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C (clk), .D (plaintext_s1[101]), .Q (new_AGEMA_signal_18901) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C (clk), .D (plaintext_s2[101]), .Q (new_AGEMA_signal_18905) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C (clk), .D (plaintext_s0[102]), .Q (new_AGEMA_signal_18909) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C (clk), .D (plaintext_s1[102]), .Q (new_AGEMA_signal_18913) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C (clk), .D (plaintext_s2[102]), .Q (new_AGEMA_signal_18917) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C (clk), .D (plaintext_s0[103]), .Q (new_AGEMA_signal_18921) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C (clk), .D (plaintext_s1[103]), .Q (new_AGEMA_signal_18925) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C (clk), .D (plaintext_s2[103]), .Q (new_AGEMA_signal_18929) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C (clk), .D (plaintext_s0[104]), .Q (new_AGEMA_signal_18933) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C (clk), .D (plaintext_s1[104]), .Q (new_AGEMA_signal_18937) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C (clk), .D (plaintext_s2[104]), .Q (new_AGEMA_signal_18941) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C (clk), .D (plaintext_s0[105]), .Q (new_AGEMA_signal_18945) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C (clk), .D (plaintext_s1[105]), .Q (new_AGEMA_signal_18949) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C (clk), .D (plaintext_s2[105]), .Q (new_AGEMA_signal_18953) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C (clk), .D (plaintext_s0[106]), .Q (new_AGEMA_signal_18957) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C (clk), .D (plaintext_s1[106]), .Q (new_AGEMA_signal_18961) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C (clk), .D (plaintext_s2[106]), .Q (new_AGEMA_signal_18965) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C (clk), .D (plaintext_s0[107]), .Q (new_AGEMA_signal_18969) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C (clk), .D (plaintext_s1[107]), .Q (new_AGEMA_signal_18973) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C (clk), .D (plaintext_s2[107]), .Q (new_AGEMA_signal_18977) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C (clk), .D (plaintext_s0[108]), .Q (new_AGEMA_signal_18981) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C (clk), .D (plaintext_s1[108]), .Q (new_AGEMA_signal_18985) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C (clk), .D (plaintext_s2[108]), .Q (new_AGEMA_signal_18989) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C (clk), .D (plaintext_s0[109]), .Q (new_AGEMA_signal_18993) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C (clk), .D (plaintext_s1[109]), .Q (new_AGEMA_signal_18997) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C (clk), .D (plaintext_s2[109]), .Q (new_AGEMA_signal_19001) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C (clk), .D (plaintext_s0[110]), .Q (new_AGEMA_signal_19005) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C (clk), .D (plaintext_s1[110]), .Q (new_AGEMA_signal_19009) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C (clk), .D (plaintext_s2[110]), .Q (new_AGEMA_signal_19013) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C (clk), .D (plaintext_s0[111]), .Q (new_AGEMA_signal_19017) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C (clk), .D (plaintext_s1[111]), .Q (new_AGEMA_signal_19021) ) ;
    buf_clk new_AGEMA_reg_buffer_6301 ( .C (clk), .D (plaintext_s2[111]), .Q (new_AGEMA_signal_19025) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C (clk), .D (plaintext_s0[112]), .Q (new_AGEMA_signal_19029) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C (clk), .D (plaintext_s1[112]), .Q (new_AGEMA_signal_19033) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C (clk), .D (plaintext_s2[112]), .Q (new_AGEMA_signal_19037) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C (clk), .D (plaintext_s0[113]), .Q (new_AGEMA_signal_19041) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C (clk), .D (plaintext_s1[113]), .Q (new_AGEMA_signal_19045) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C (clk), .D (plaintext_s2[113]), .Q (new_AGEMA_signal_19049) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C (clk), .D (plaintext_s0[114]), .Q (new_AGEMA_signal_19053) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C (clk), .D (plaintext_s1[114]), .Q (new_AGEMA_signal_19057) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C (clk), .D (plaintext_s2[114]), .Q (new_AGEMA_signal_19061) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C (clk), .D (plaintext_s0[115]), .Q (new_AGEMA_signal_19065) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C (clk), .D (plaintext_s1[115]), .Q (new_AGEMA_signal_19069) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C (clk), .D (plaintext_s2[115]), .Q (new_AGEMA_signal_19073) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C (clk), .D (plaintext_s0[116]), .Q (new_AGEMA_signal_19077) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C (clk), .D (plaintext_s1[116]), .Q (new_AGEMA_signal_19081) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C (clk), .D (plaintext_s2[116]), .Q (new_AGEMA_signal_19085) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C (clk), .D (plaintext_s0[117]), .Q (new_AGEMA_signal_19089) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C (clk), .D (plaintext_s1[117]), .Q (new_AGEMA_signal_19093) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C (clk), .D (plaintext_s2[117]), .Q (new_AGEMA_signal_19097) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C (clk), .D (plaintext_s0[118]), .Q (new_AGEMA_signal_19101) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C (clk), .D (plaintext_s1[118]), .Q (new_AGEMA_signal_19105) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C (clk), .D (plaintext_s2[118]), .Q (new_AGEMA_signal_19109) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C (clk), .D (plaintext_s0[119]), .Q (new_AGEMA_signal_19113) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C (clk), .D (plaintext_s1[119]), .Q (new_AGEMA_signal_19117) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C (clk), .D (plaintext_s2[119]), .Q (new_AGEMA_signal_19121) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C (clk), .D (plaintext_s0[120]), .Q (new_AGEMA_signal_19125) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C (clk), .D (plaintext_s1[120]), .Q (new_AGEMA_signal_19129) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C (clk), .D (plaintext_s2[120]), .Q (new_AGEMA_signal_19133) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C (clk), .D (plaintext_s0[121]), .Q (new_AGEMA_signal_19137) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C (clk), .D (plaintext_s1[121]), .Q (new_AGEMA_signal_19141) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C (clk), .D (plaintext_s2[121]), .Q (new_AGEMA_signal_19145) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C (clk), .D (plaintext_s0[122]), .Q (new_AGEMA_signal_19149) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C (clk), .D (plaintext_s1[122]), .Q (new_AGEMA_signal_19153) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C (clk), .D (plaintext_s2[122]), .Q (new_AGEMA_signal_19157) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C (clk), .D (plaintext_s0[123]), .Q (new_AGEMA_signal_19161) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C (clk), .D (plaintext_s1[123]), .Q (new_AGEMA_signal_19165) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C (clk), .D (plaintext_s2[123]), .Q (new_AGEMA_signal_19169) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C (clk), .D (plaintext_s0[124]), .Q (new_AGEMA_signal_19173) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C (clk), .D (plaintext_s1[124]), .Q (new_AGEMA_signal_19177) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C (clk), .D (plaintext_s2[124]), .Q (new_AGEMA_signal_19181) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C (clk), .D (plaintext_s0[125]), .Q (new_AGEMA_signal_19185) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C (clk), .D (plaintext_s1[125]), .Q (new_AGEMA_signal_19189) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C (clk), .D (plaintext_s2[125]), .Q (new_AGEMA_signal_19193) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C (clk), .D (plaintext_s0[126]), .Q (new_AGEMA_signal_19197) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C (clk), .D (plaintext_s1[126]), .Q (new_AGEMA_signal_19201) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C (clk), .D (plaintext_s2[126]), .Q (new_AGEMA_signal_19205) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C (clk), .D (plaintext_s0[127]), .Q (new_AGEMA_signal_19209) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C (clk), .D (plaintext_s1[127]), .Q (new_AGEMA_signal_19213) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C (clk), .D (plaintext_s2[127]), .Q (new_AGEMA_signal_19217) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_19221) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_5781), .Q (new_AGEMA_signal_19224) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_19227) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_19230) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C (clk), .D (new_AGEMA_signal_6141), .Q (new_AGEMA_signal_19233) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_19236) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_19239) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_19242) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C (clk), .D (ciphertext_s2[0]), .Q (new_AGEMA_signal_19245) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_19248) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_5789), .Q (new_AGEMA_signal_19251) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_19254) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_19257) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_19260) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_19263) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_19266) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_19269) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_19272) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_19275) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_19278) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_19281) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_19284) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_19287) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_19290) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_19293) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_19296) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_19299) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_19302) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C (clk), .D (new_AGEMA_signal_5785), .Q (new_AGEMA_signal_19305) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_19308) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_19311) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_19314) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_19317) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_19320) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_19323) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_19326) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_19329) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_19332) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_19335) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_19338) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_19341) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_19344) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_19347) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_6149), .Q (new_AGEMA_signal_19350) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_19353) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_19356) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_19359) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_19362) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_19365) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_19368) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_19371) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_19374) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_19377) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_19380) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_19383) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_5797), .Q (new_AGEMA_signal_19386) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_19389) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_19392) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_19395) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_19398) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_19401) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_19404) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C (clk), .D (ciphertext_s2[8]), .Q (new_AGEMA_signal_19407) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_19410) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C (clk), .D (new_AGEMA_signal_5805), .Q (new_AGEMA_signal_19413) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_19416) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_19419) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_19422) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_19425) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_19428) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C (clk), .D (new_AGEMA_signal_6173), .Q (new_AGEMA_signal_19431) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_19434) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_19437) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_19440) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_19443) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_19446) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_19449) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_19452) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_19455) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C (clk), .D (new_AGEMA_signal_6169), .Q (new_AGEMA_signal_19458) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_19461) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_19464) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_19467) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_19470) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_19473) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_19476) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C (clk), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_19479) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_19482) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_19485) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_19488) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_19491) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C (clk), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_19494) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C (clk), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_19497) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_19500) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C (clk), .D (new_AGEMA_signal_5809), .Q (new_AGEMA_signal_19503) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_19506) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_19509) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_19512) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_19515) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_19518) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C (clk), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_19521) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_19524) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_19527) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_19530) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_19533) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_19536) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_19539) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_19542) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_19545) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C (clk), .D (new_AGEMA_signal_5813), .Q (new_AGEMA_signal_19548) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_19551) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_19554) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C (clk), .D (new_AGEMA_signal_6193), .Q (new_AGEMA_signal_19557) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_19560) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_19563) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_19566) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C (clk), .D (ciphertext_s2[16]), .Q (new_AGEMA_signal_19569) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_19572) ) ;
    buf_clk new_AGEMA_reg_buffer_6851 ( .C (clk), .D (new_AGEMA_signal_5821), .Q (new_AGEMA_signal_19575) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_19578) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_19581) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_19584) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_19587) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_19590) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_19593) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_19596) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_19599) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_19602) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_19605) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_19608) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_19611) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_19614) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_19617) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_19620) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_19623) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_19626) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_19629) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C (clk), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_19632) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_19635) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_19638) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_19641) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_19644) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_19647) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_19650) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_19653) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C (clk), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_19656) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_19659) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_19662) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_19665) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_19668) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_19671) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_19674) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C (clk), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_19677) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_19680) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_19683) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_19686) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_19689) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_19692) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_19695) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_19698) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_19701) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_19704) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_19707) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_19710) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_19713) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_19716) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_19719) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_19722) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_19725) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_19728) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C (clk), .D (ciphertext_s2[24]), .Q (new_AGEMA_signal_19731) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_19734) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C (clk), .D (new_AGEMA_signal_5837), .Q (new_AGEMA_signal_19737) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_19740) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_19743) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_19746) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_19749) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_19752) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_19755) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C (clk), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_19758) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_19761) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_19764) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_19767) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_19770) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_19773) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_19776) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_19779) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C (clk), .D (new_AGEMA_signal_6221), .Q (new_AGEMA_signal_19782) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_19785) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_19788) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C (clk), .D (new_AGEMA_signal_5833), .Q (new_AGEMA_signal_19791) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_19794) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_19797) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C (clk), .D (new_AGEMA_signal_6229), .Q (new_AGEMA_signal_19800) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_19803) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_19806) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_19809) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_19812) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_19815) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_19818) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_19821) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_19824) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_19827) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C (clk), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_19830) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_19833) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_19836) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_19839) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_19842) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C (clk), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_19845) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C (clk), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_19848) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_19851) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_19854) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_19857) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_19860) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C (clk), .D (new_AGEMA_signal_5459), .Q (new_AGEMA_signal_19863) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_19866) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T6), .Q (new_AGEMA_signal_19869) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C (clk), .D (new_AGEMA_signal_5845), .Q (new_AGEMA_signal_19872) ) ;
    buf_clk new_AGEMA_reg_buffer_7151 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_19875) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T8), .Q (new_AGEMA_signal_19878) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C (clk), .D (new_AGEMA_signal_6245), .Q (new_AGEMA_signal_19881) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_19884) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_19887) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_19890) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C (clk), .D (ciphertext_s2[32]), .Q (new_AGEMA_signal_19893) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T16), .Q (new_AGEMA_signal_19896) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_19899) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_19902) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T9), .Q (new_AGEMA_signal_19905) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_19908) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_19911) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T17), .Q (new_AGEMA_signal_19914) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_19917) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_19920) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T15), .Q (new_AGEMA_signal_19923) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_19926) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_19929) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T27), .Q (new_AGEMA_signal_19932) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_19935) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_19938) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T10), .Q (new_AGEMA_signal_19941) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_19944) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_19947) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T13), .Q (new_AGEMA_signal_19950) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C (clk), .D (new_AGEMA_signal_5849), .Q (new_AGEMA_signal_19953) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_19956) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T23), .Q (new_AGEMA_signal_19959) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_19962) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_19965) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T19), .Q (new_AGEMA_signal_19968) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_19971) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_19974) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T3), .Q (new_AGEMA_signal_19977) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_19980) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C (clk), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_19983) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T22), .Q (new_AGEMA_signal_19986) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_19989) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_19992) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T20), .Q (new_AGEMA_signal_19995) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C (clk), .D (new_AGEMA_signal_6253), .Q (new_AGEMA_signal_19998) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_20001) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T1), .Q (new_AGEMA_signal_20004) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C (clk), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_20007) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_20010) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T4), .Q (new_AGEMA_signal_20013) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C (clk), .D (new_AGEMA_signal_5483), .Q (new_AGEMA_signal_20016) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_20019) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_T2), .Q (new_AGEMA_signal_20022) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_20025) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_20028) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T6), .Q (new_AGEMA_signal_20031) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C (clk), .D (new_AGEMA_signal_5861), .Q (new_AGEMA_signal_20034) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_20037) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T8), .Q (new_AGEMA_signal_20040) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_20043) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_20046) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_20049) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_20052) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C (clk), .D (ciphertext_s2[40]), .Q (new_AGEMA_signal_20055) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T16), .Q (new_AGEMA_signal_20058) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C (clk), .D (new_AGEMA_signal_5869), .Q (new_AGEMA_signal_20061) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_20064) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T9), .Q (new_AGEMA_signal_20067) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_20070) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_20073) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T17), .Q (new_AGEMA_signal_20076) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C (clk), .D (new_AGEMA_signal_6277), .Q (new_AGEMA_signal_20079) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_20082) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T15), .Q (new_AGEMA_signal_20085) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_20088) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_20091) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T27), .Q (new_AGEMA_signal_20094) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_20097) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_20100) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T10), .Q (new_AGEMA_signal_20103) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_20106) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_20109) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T13), .Q (new_AGEMA_signal_20112) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_20115) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C (clk), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_20118) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T23), .Q (new_AGEMA_signal_20121) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C (clk), .D (new_AGEMA_signal_6281), .Q (new_AGEMA_signal_20124) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_20127) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T19), .Q (new_AGEMA_signal_20130) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_20133) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_20136) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T3), .Q (new_AGEMA_signal_20139) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_20142) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_20145) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T22), .Q (new_AGEMA_signal_20148) ) ;
    buf_clk new_AGEMA_reg_buffer_7427 ( .C (clk), .D (new_AGEMA_signal_5873), .Q (new_AGEMA_signal_20151) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_20154) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T20), .Q (new_AGEMA_signal_20157) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_20160) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_20163) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T1), .Q (new_AGEMA_signal_20166) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_20169) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_20172) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T4), .Q (new_AGEMA_signal_20175) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_20178) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_20181) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_T2), .Q (new_AGEMA_signal_20184) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_20187) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_20190) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T6), .Q (new_AGEMA_signal_20193) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C (clk), .D (new_AGEMA_signal_5877), .Q (new_AGEMA_signal_20196) ) ;
    buf_clk new_AGEMA_reg_buffer_7475 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_20199) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T8), .Q (new_AGEMA_signal_20202) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C (clk), .D (new_AGEMA_signal_6297), .Q (new_AGEMA_signal_20205) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C (clk), .D (new_AGEMA_signal_6298), .Q (new_AGEMA_signal_20208) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_20211) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_20214) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C (clk), .D (ciphertext_s2[48]), .Q (new_AGEMA_signal_20217) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T16), .Q (new_AGEMA_signal_20220) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C (clk), .D (new_AGEMA_signal_5885), .Q (new_AGEMA_signal_20223) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_20226) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T9), .Q (new_AGEMA_signal_20229) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_20232) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_20235) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T17), .Q (new_AGEMA_signal_20238) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_20241) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_20244) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T15), .Q (new_AGEMA_signal_20247) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_20250) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_20253) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T27), .Q (new_AGEMA_signal_20256) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_20259) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_20262) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T10), .Q (new_AGEMA_signal_20265) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_20268) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_20271) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T13), .Q (new_AGEMA_signal_20274) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_20277) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_20280) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T23), .Q (new_AGEMA_signal_20283) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_20286) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_20289) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T19), .Q (new_AGEMA_signal_20292) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_20295) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_20298) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T3), .Q (new_AGEMA_signal_20301) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_20304) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_20307) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T22), .Q (new_AGEMA_signal_20310) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_20313) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_20316) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T20), .Q (new_AGEMA_signal_20319) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C (clk), .D (new_AGEMA_signal_6305), .Q (new_AGEMA_signal_20322) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_20325) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T1), .Q (new_AGEMA_signal_20328) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_20331) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_20334) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T4), .Q (new_AGEMA_signal_20337) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_20340) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_20343) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_T2), .Q (new_AGEMA_signal_20346) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_20349) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_20352) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T6), .Q (new_AGEMA_signal_20355) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C (clk), .D (new_AGEMA_signal_5893), .Q (new_AGEMA_signal_20358) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_20361) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T8), .Q (new_AGEMA_signal_20364) ) ;
    buf_clk new_AGEMA_reg_buffer_7643 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_20367) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_20370) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_20373) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_20376) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C (clk), .D (ciphertext_s2[56]), .Q (new_AGEMA_signal_20379) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T16), .Q (new_AGEMA_signal_20382) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C (clk), .D (new_AGEMA_signal_5901), .Q (new_AGEMA_signal_20385) ) ;
    buf_clk new_AGEMA_reg_buffer_7664 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_20388) ) ;
    buf_clk new_AGEMA_reg_buffer_7667 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T9), .Q (new_AGEMA_signal_20391) ) ;
    buf_clk new_AGEMA_reg_buffer_7670 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_20394) ) ;
    buf_clk new_AGEMA_reg_buffer_7673 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_20397) ) ;
    buf_clk new_AGEMA_reg_buffer_7676 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T17), .Q (new_AGEMA_signal_20400) ) ;
    buf_clk new_AGEMA_reg_buffer_7679 ( .C (clk), .D (new_AGEMA_signal_6329), .Q (new_AGEMA_signal_20403) ) ;
    buf_clk new_AGEMA_reg_buffer_7682 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_20406) ) ;
    buf_clk new_AGEMA_reg_buffer_7685 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T15), .Q (new_AGEMA_signal_20409) ) ;
    buf_clk new_AGEMA_reg_buffer_7688 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_20412) ) ;
    buf_clk new_AGEMA_reg_buffer_7691 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_20415) ) ;
    buf_clk new_AGEMA_reg_buffer_7694 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T27), .Q (new_AGEMA_signal_20418) ) ;
    buf_clk new_AGEMA_reg_buffer_7697 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_20421) ) ;
    buf_clk new_AGEMA_reg_buffer_7700 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_20424) ) ;
    buf_clk new_AGEMA_reg_buffer_7703 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T10), .Q (new_AGEMA_signal_20427) ) ;
    buf_clk new_AGEMA_reg_buffer_7706 ( .C (clk), .D (new_AGEMA_signal_6325), .Q (new_AGEMA_signal_20430) ) ;
    buf_clk new_AGEMA_reg_buffer_7709 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_20433) ) ;
    buf_clk new_AGEMA_reg_buffer_7712 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T13), .Q (new_AGEMA_signal_20436) ) ;
    buf_clk new_AGEMA_reg_buffer_7715 ( .C (clk), .D (new_AGEMA_signal_5897), .Q (new_AGEMA_signal_20439) ) ;
    buf_clk new_AGEMA_reg_buffer_7718 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_20442) ) ;
    buf_clk new_AGEMA_reg_buffer_7721 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T23), .Q (new_AGEMA_signal_20445) ) ;
    buf_clk new_AGEMA_reg_buffer_7724 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_20448) ) ;
    buf_clk new_AGEMA_reg_buffer_7727 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_20451) ) ;
    buf_clk new_AGEMA_reg_buffer_7730 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T19), .Q (new_AGEMA_signal_20454) ) ;
    buf_clk new_AGEMA_reg_buffer_7733 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_20457) ) ;
    buf_clk new_AGEMA_reg_buffer_7736 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_20460) ) ;
    buf_clk new_AGEMA_reg_buffer_7739 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T3), .Q (new_AGEMA_signal_20463) ) ;
    buf_clk new_AGEMA_reg_buffer_7742 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_20466) ) ;
    buf_clk new_AGEMA_reg_buffer_7745 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_20469) ) ;
    buf_clk new_AGEMA_reg_buffer_7748 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T22), .Q (new_AGEMA_signal_20472) ) ;
    buf_clk new_AGEMA_reg_buffer_7751 ( .C (clk), .D (new_AGEMA_signal_5905), .Q (new_AGEMA_signal_20475) ) ;
    buf_clk new_AGEMA_reg_buffer_7754 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_20478) ) ;
    buf_clk new_AGEMA_reg_buffer_7757 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T20), .Q (new_AGEMA_signal_20481) ) ;
    buf_clk new_AGEMA_reg_buffer_7760 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_20484) ) ;
    buf_clk new_AGEMA_reg_buffer_7763 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_20487) ) ;
    buf_clk new_AGEMA_reg_buffer_7766 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T1), .Q (new_AGEMA_signal_20490) ) ;
    buf_clk new_AGEMA_reg_buffer_7769 ( .C (clk), .D (new_AGEMA_signal_5537), .Q (new_AGEMA_signal_20493) ) ;
    buf_clk new_AGEMA_reg_buffer_7772 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_20496) ) ;
    buf_clk new_AGEMA_reg_buffer_7775 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T4), .Q (new_AGEMA_signal_20499) ) ;
    buf_clk new_AGEMA_reg_buffer_7778 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_20502) ) ;
    buf_clk new_AGEMA_reg_buffer_7781 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_20505) ) ;
    buf_clk new_AGEMA_reg_buffer_7784 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_T2), .Q (new_AGEMA_signal_20508) ) ;
    buf_clk new_AGEMA_reg_buffer_7787 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_20511) ) ;
    buf_clk new_AGEMA_reg_buffer_7790 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_20514) ) ;
    buf_clk new_AGEMA_reg_buffer_7793 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T6), .Q (new_AGEMA_signal_20517) ) ;
    buf_clk new_AGEMA_reg_buffer_7796 ( .C (clk), .D (new_AGEMA_signal_5909), .Q (new_AGEMA_signal_20520) ) ;
    buf_clk new_AGEMA_reg_buffer_7799 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_20523) ) ;
    buf_clk new_AGEMA_reg_buffer_7802 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T8), .Q (new_AGEMA_signal_20526) ) ;
    buf_clk new_AGEMA_reg_buffer_7805 ( .C (clk), .D (new_AGEMA_signal_6349), .Q (new_AGEMA_signal_20529) ) ;
    buf_clk new_AGEMA_reg_buffer_7808 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_20532) ) ;
    buf_clk new_AGEMA_reg_buffer_7811 ( .C (clk), .D (ciphertext_s0[64]), .Q (new_AGEMA_signal_20535) ) ;
    buf_clk new_AGEMA_reg_buffer_7814 ( .C (clk), .D (ciphertext_s1[64]), .Q (new_AGEMA_signal_20538) ) ;
    buf_clk new_AGEMA_reg_buffer_7817 ( .C (clk), .D (ciphertext_s2[64]), .Q (new_AGEMA_signal_20541) ) ;
    buf_clk new_AGEMA_reg_buffer_7820 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T16), .Q (new_AGEMA_signal_20544) ) ;
    buf_clk new_AGEMA_reg_buffer_7823 ( .C (clk), .D (new_AGEMA_signal_5917), .Q (new_AGEMA_signal_20547) ) ;
    buf_clk new_AGEMA_reg_buffer_7826 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_20550) ) ;
    buf_clk new_AGEMA_reg_buffer_7829 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T9), .Q (new_AGEMA_signal_20553) ) ;
    buf_clk new_AGEMA_reg_buffer_7832 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_20556) ) ;
    buf_clk new_AGEMA_reg_buffer_7835 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_20559) ) ;
    buf_clk new_AGEMA_reg_buffer_7838 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T17), .Q (new_AGEMA_signal_20562) ) ;
    buf_clk new_AGEMA_reg_buffer_7841 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_20565) ) ;
    buf_clk new_AGEMA_reg_buffer_7844 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_20568) ) ;
    buf_clk new_AGEMA_reg_buffer_7847 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T15), .Q (new_AGEMA_signal_20571) ) ;
    buf_clk new_AGEMA_reg_buffer_7850 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_20574) ) ;
    buf_clk new_AGEMA_reg_buffer_7853 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_20577) ) ;
    buf_clk new_AGEMA_reg_buffer_7856 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T27), .Q (new_AGEMA_signal_20580) ) ;
    buf_clk new_AGEMA_reg_buffer_7859 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_20583) ) ;
    buf_clk new_AGEMA_reg_buffer_7862 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_20586) ) ;
    buf_clk new_AGEMA_reg_buffer_7865 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T10), .Q (new_AGEMA_signal_20589) ) ;
    buf_clk new_AGEMA_reg_buffer_7868 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_20592) ) ;
    buf_clk new_AGEMA_reg_buffer_7871 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_20595) ) ;
    buf_clk new_AGEMA_reg_buffer_7874 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T13), .Q (new_AGEMA_signal_20598) ) ;
    buf_clk new_AGEMA_reg_buffer_7877 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_20601) ) ;
    buf_clk new_AGEMA_reg_buffer_7880 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_20604) ) ;
    buf_clk new_AGEMA_reg_buffer_7883 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T23), .Q (new_AGEMA_signal_20607) ) ;
    buf_clk new_AGEMA_reg_buffer_7886 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_20610) ) ;
    buf_clk new_AGEMA_reg_buffer_7889 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_20613) ) ;
    buf_clk new_AGEMA_reg_buffer_7892 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T19), .Q (new_AGEMA_signal_20616) ) ;
    buf_clk new_AGEMA_reg_buffer_7895 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_20619) ) ;
    buf_clk new_AGEMA_reg_buffer_7898 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_20622) ) ;
    buf_clk new_AGEMA_reg_buffer_7901 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T3), .Q (new_AGEMA_signal_20625) ) ;
    buf_clk new_AGEMA_reg_buffer_7904 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_20628) ) ;
    buf_clk new_AGEMA_reg_buffer_7907 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_20631) ) ;
    buf_clk new_AGEMA_reg_buffer_7910 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T22), .Q (new_AGEMA_signal_20634) ) ;
    buf_clk new_AGEMA_reg_buffer_7913 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_20637) ) ;
    buf_clk new_AGEMA_reg_buffer_7916 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_20640) ) ;
    buf_clk new_AGEMA_reg_buffer_7919 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T20), .Q (new_AGEMA_signal_20643) ) ;
    buf_clk new_AGEMA_reg_buffer_7922 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_20646) ) ;
    buf_clk new_AGEMA_reg_buffer_7925 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_20649) ) ;
    buf_clk new_AGEMA_reg_buffer_7928 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T1), .Q (new_AGEMA_signal_20652) ) ;
    buf_clk new_AGEMA_reg_buffer_7931 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_20655) ) ;
    buf_clk new_AGEMA_reg_buffer_7934 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_20658) ) ;
    buf_clk new_AGEMA_reg_buffer_7937 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T4), .Q (new_AGEMA_signal_20661) ) ;
    buf_clk new_AGEMA_reg_buffer_7940 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_20664) ) ;
    buf_clk new_AGEMA_reg_buffer_7943 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_20667) ) ;
    buf_clk new_AGEMA_reg_buffer_7946 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_T2), .Q (new_AGEMA_signal_20670) ) ;
    buf_clk new_AGEMA_reg_buffer_7949 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_20673) ) ;
    buf_clk new_AGEMA_reg_buffer_7952 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_20676) ) ;
    buf_clk new_AGEMA_reg_buffer_7955 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T6), .Q (new_AGEMA_signal_20679) ) ;
    buf_clk new_AGEMA_reg_buffer_7958 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_20682) ) ;
    buf_clk new_AGEMA_reg_buffer_7961 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_20685) ) ;
    buf_clk new_AGEMA_reg_buffer_7964 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T8), .Q (new_AGEMA_signal_20688) ) ;
    buf_clk new_AGEMA_reg_buffer_7967 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_20691) ) ;
    buf_clk new_AGEMA_reg_buffer_7970 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_20694) ) ;
    buf_clk new_AGEMA_reg_buffer_7973 ( .C (clk), .D (ciphertext_s0[72]), .Q (new_AGEMA_signal_20697) ) ;
    buf_clk new_AGEMA_reg_buffer_7976 ( .C (clk), .D (ciphertext_s1[72]), .Q (new_AGEMA_signal_20700) ) ;
    buf_clk new_AGEMA_reg_buffer_7979 ( .C (clk), .D (ciphertext_s2[72]), .Q (new_AGEMA_signal_20703) ) ;
    buf_clk new_AGEMA_reg_buffer_7982 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T16), .Q (new_AGEMA_signal_20706) ) ;
    buf_clk new_AGEMA_reg_buffer_7985 ( .C (clk), .D (new_AGEMA_signal_5933), .Q (new_AGEMA_signal_20709) ) ;
    buf_clk new_AGEMA_reg_buffer_7988 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_20712) ) ;
    buf_clk new_AGEMA_reg_buffer_7991 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T9), .Q (new_AGEMA_signal_20715) ) ;
    buf_clk new_AGEMA_reg_buffer_7994 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_20718) ) ;
    buf_clk new_AGEMA_reg_buffer_7997 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_20721) ) ;
    buf_clk new_AGEMA_reg_buffer_8000 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T17), .Q (new_AGEMA_signal_20724) ) ;
    buf_clk new_AGEMA_reg_buffer_8003 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_20727) ) ;
    buf_clk new_AGEMA_reg_buffer_8006 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_20730) ) ;
    buf_clk new_AGEMA_reg_buffer_8009 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T15), .Q (new_AGEMA_signal_20733) ) ;
    buf_clk new_AGEMA_reg_buffer_8012 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_20736) ) ;
    buf_clk new_AGEMA_reg_buffer_8015 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_20739) ) ;
    buf_clk new_AGEMA_reg_buffer_8018 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T27), .Q (new_AGEMA_signal_20742) ) ;
    buf_clk new_AGEMA_reg_buffer_8021 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_20745) ) ;
    buf_clk new_AGEMA_reg_buffer_8024 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_20748) ) ;
    buf_clk new_AGEMA_reg_buffer_8027 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T10), .Q (new_AGEMA_signal_20751) ) ;
    buf_clk new_AGEMA_reg_buffer_8030 ( .C (clk), .D (new_AGEMA_signal_6377), .Q (new_AGEMA_signal_20754) ) ;
    buf_clk new_AGEMA_reg_buffer_8033 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_20757) ) ;
    buf_clk new_AGEMA_reg_buffer_8036 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T13), .Q (new_AGEMA_signal_20760) ) ;
    buf_clk new_AGEMA_reg_buffer_8039 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_20763) ) ;
    buf_clk new_AGEMA_reg_buffer_8042 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_20766) ) ;
    buf_clk new_AGEMA_reg_buffer_8045 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T23), .Q (new_AGEMA_signal_20769) ) ;
    buf_clk new_AGEMA_reg_buffer_8048 ( .C (clk), .D (new_AGEMA_signal_6385), .Q (new_AGEMA_signal_20772) ) ;
    buf_clk new_AGEMA_reg_buffer_8051 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_20775) ) ;
    buf_clk new_AGEMA_reg_buffer_8054 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T19), .Q (new_AGEMA_signal_20778) ) ;
    buf_clk new_AGEMA_reg_buffer_8057 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_20781) ) ;
    buf_clk new_AGEMA_reg_buffer_8060 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_20784) ) ;
    buf_clk new_AGEMA_reg_buffer_8063 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T3), .Q (new_AGEMA_signal_20787) ) ;
    buf_clk new_AGEMA_reg_buffer_8066 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_20790) ) ;
    buf_clk new_AGEMA_reg_buffer_8069 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_20793) ) ;
    buf_clk new_AGEMA_reg_buffer_8072 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T22), .Q (new_AGEMA_signal_20796) ) ;
    buf_clk new_AGEMA_reg_buffer_8075 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_20799) ) ;
    buf_clk new_AGEMA_reg_buffer_8078 ( .C (clk), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_20802) ) ;
    buf_clk new_AGEMA_reg_buffer_8081 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T20), .Q (new_AGEMA_signal_20805) ) ;
    buf_clk new_AGEMA_reg_buffer_8084 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_20808) ) ;
    buf_clk new_AGEMA_reg_buffer_8087 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_20811) ) ;
    buf_clk new_AGEMA_reg_buffer_8090 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T1), .Q (new_AGEMA_signal_20814) ) ;
    buf_clk new_AGEMA_reg_buffer_8093 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_20817) ) ;
    buf_clk new_AGEMA_reg_buffer_8096 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_20820) ) ;
    buf_clk new_AGEMA_reg_buffer_8099 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T4), .Q (new_AGEMA_signal_20823) ) ;
    buf_clk new_AGEMA_reg_buffer_8102 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_20826) ) ;
    buf_clk new_AGEMA_reg_buffer_8105 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_20829) ) ;
    buf_clk new_AGEMA_reg_buffer_8108 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_T2), .Q (new_AGEMA_signal_20832) ) ;
    buf_clk new_AGEMA_reg_buffer_8111 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_20835) ) ;
    buf_clk new_AGEMA_reg_buffer_8114 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_20838) ) ;
    buf_clk new_AGEMA_reg_buffer_8117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T6), .Q (new_AGEMA_signal_20841) ) ;
    buf_clk new_AGEMA_reg_buffer_8120 ( .C (clk), .D (new_AGEMA_signal_5941), .Q (new_AGEMA_signal_20844) ) ;
    buf_clk new_AGEMA_reg_buffer_8123 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_20847) ) ;
    buf_clk new_AGEMA_reg_buffer_8126 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T8), .Q (new_AGEMA_signal_20850) ) ;
    buf_clk new_AGEMA_reg_buffer_8129 ( .C (clk), .D (new_AGEMA_signal_6401), .Q (new_AGEMA_signal_20853) ) ;
    buf_clk new_AGEMA_reg_buffer_8132 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_20856) ) ;
    buf_clk new_AGEMA_reg_buffer_8135 ( .C (clk), .D (ciphertext_s0[80]), .Q (new_AGEMA_signal_20859) ) ;
    buf_clk new_AGEMA_reg_buffer_8138 ( .C (clk), .D (ciphertext_s1[80]), .Q (new_AGEMA_signal_20862) ) ;
    buf_clk new_AGEMA_reg_buffer_8141 ( .C (clk), .D (ciphertext_s2[80]), .Q (new_AGEMA_signal_20865) ) ;
    buf_clk new_AGEMA_reg_buffer_8144 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T16), .Q (new_AGEMA_signal_20868) ) ;
    buf_clk new_AGEMA_reg_buffer_8147 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_20871) ) ;
    buf_clk new_AGEMA_reg_buffer_8150 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_20874) ) ;
    buf_clk new_AGEMA_reg_buffer_8153 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T9), .Q (new_AGEMA_signal_20877) ) ;
    buf_clk new_AGEMA_reg_buffer_8156 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_20880) ) ;
    buf_clk new_AGEMA_reg_buffer_8159 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_20883) ) ;
    buf_clk new_AGEMA_reg_buffer_8162 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T17), .Q (new_AGEMA_signal_20886) ) ;
    buf_clk new_AGEMA_reg_buffer_8165 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_20889) ) ;
    buf_clk new_AGEMA_reg_buffer_8168 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_20892) ) ;
    buf_clk new_AGEMA_reg_buffer_8171 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T15), .Q (new_AGEMA_signal_20895) ) ;
    buf_clk new_AGEMA_reg_buffer_8174 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_20898) ) ;
    buf_clk new_AGEMA_reg_buffer_8177 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_20901) ) ;
    buf_clk new_AGEMA_reg_buffer_8180 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T27), .Q (new_AGEMA_signal_20904) ) ;
    buf_clk new_AGEMA_reg_buffer_8183 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_20907) ) ;
    buf_clk new_AGEMA_reg_buffer_8186 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_20910) ) ;
    buf_clk new_AGEMA_reg_buffer_8189 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T10), .Q (new_AGEMA_signal_20913) ) ;
    buf_clk new_AGEMA_reg_buffer_8192 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_20916) ) ;
    buf_clk new_AGEMA_reg_buffer_8195 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_20919) ) ;
    buf_clk new_AGEMA_reg_buffer_8198 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T13), .Q (new_AGEMA_signal_20922) ) ;
    buf_clk new_AGEMA_reg_buffer_8201 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_20925) ) ;
    buf_clk new_AGEMA_reg_buffer_8204 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_20928) ) ;
    buf_clk new_AGEMA_reg_buffer_8207 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T23), .Q (new_AGEMA_signal_20931) ) ;
    buf_clk new_AGEMA_reg_buffer_8210 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_20934) ) ;
    buf_clk new_AGEMA_reg_buffer_8213 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_20937) ) ;
    buf_clk new_AGEMA_reg_buffer_8216 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T19), .Q (new_AGEMA_signal_20940) ) ;
    buf_clk new_AGEMA_reg_buffer_8219 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_20943) ) ;
    buf_clk new_AGEMA_reg_buffer_8222 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_20946) ) ;
    buf_clk new_AGEMA_reg_buffer_8225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T3), .Q (new_AGEMA_signal_20949) ) ;
    buf_clk new_AGEMA_reg_buffer_8228 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_20952) ) ;
    buf_clk new_AGEMA_reg_buffer_8231 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_20955) ) ;
    buf_clk new_AGEMA_reg_buffer_8234 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T22), .Q (new_AGEMA_signal_20958) ) ;
    buf_clk new_AGEMA_reg_buffer_8237 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_20961) ) ;
    buf_clk new_AGEMA_reg_buffer_8240 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_20964) ) ;
    buf_clk new_AGEMA_reg_buffer_8243 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T20), .Q (new_AGEMA_signal_20967) ) ;
    buf_clk new_AGEMA_reg_buffer_8246 ( .C (clk), .D (new_AGEMA_signal_6409), .Q (new_AGEMA_signal_20970) ) ;
    buf_clk new_AGEMA_reg_buffer_8249 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_20973) ) ;
    buf_clk new_AGEMA_reg_buffer_8252 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T1), .Q (new_AGEMA_signal_20976) ) ;
    buf_clk new_AGEMA_reg_buffer_8255 ( .C (clk), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_20979) ) ;
    buf_clk new_AGEMA_reg_buffer_8258 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_20982) ) ;
    buf_clk new_AGEMA_reg_buffer_8261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T4), .Q (new_AGEMA_signal_20985) ) ;
    buf_clk new_AGEMA_reg_buffer_8264 ( .C (clk), .D (new_AGEMA_signal_5603), .Q (new_AGEMA_signal_20988) ) ;
    buf_clk new_AGEMA_reg_buffer_8267 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_20991) ) ;
    buf_clk new_AGEMA_reg_buffer_8270 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_T2), .Q (new_AGEMA_signal_20994) ) ;
    buf_clk new_AGEMA_reg_buffer_8273 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_20997) ) ;
    buf_clk new_AGEMA_reg_buffer_8276 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_21000) ) ;
    buf_clk new_AGEMA_reg_buffer_8279 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T6), .Q (new_AGEMA_signal_21003) ) ;
    buf_clk new_AGEMA_reg_buffer_8282 ( .C (clk), .D (new_AGEMA_signal_5957), .Q (new_AGEMA_signal_21006) ) ;
    buf_clk new_AGEMA_reg_buffer_8285 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_21009) ) ;
    buf_clk new_AGEMA_reg_buffer_8288 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T8), .Q (new_AGEMA_signal_21012) ) ;
    buf_clk new_AGEMA_reg_buffer_8291 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_21015) ) ;
    buf_clk new_AGEMA_reg_buffer_8294 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_21018) ) ;
    buf_clk new_AGEMA_reg_buffer_8297 ( .C (clk), .D (ciphertext_s0[88]), .Q (new_AGEMA_signal_21021) ) ;
    buf_clk new_AGEMA_reg_buffer_8300 ( .C (clk), .D (ciphertext_s1[88]), .Q (new_AGEMA_signal_21024) ) ;
    buf_clk new_AGEMA_reg_buffer_8303 ( .C (clk), .D (ciphertext_s2[88]), .Q (new_AGEMA_signal_21027) ) ;
    buf_clk new_AGEMA_reg_buffer_8306 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T16), .Q (new_AGEMA_signal_21030) ) ;
    buf_clk new_AGEMA_reg_buffer_8309 ( .C (clk), .D (new_AGEMA_signal_5965), .Q (new_AGEMA_signal_21033) ) ;
    buf_clk new_AGEMA_reg_buffer_8312 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_21036) ) ;
    buf_clk new_AGEMA_reg_buffer_8315 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T9), .Q (new_AGEMA_signal_21039) ) ;
    buf_clk new_AGEMA_reg_buffer_8318 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_21042) ) ;
    buf_clk new_AGEMA_reg_buffer_8321 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_21045) ) ;
    buf_clk new_AGEMA_reg_buffer_8324 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T17), .Q (new_AGEMA_signal_21048) ) ;
    buf_clk new_AGEMA_reg_buffer_8327 ( .C (clk), .D (new_AGEMA_signal_6433), .Q (new_AGEMA_signal_21051) ) ;
    buf_clk new_AGEMA_reg_buffer_8330 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_21054) ) ;
    buf_clk new_AGEMA_reg_buffer_8333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T15), .Q (new_AGEMA_signal_21057) ) ;
    buf_clk new_AGEMA_reg_buffer_8336 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_21060) ) ;
    buf_clk new_AGEMA_reg_buffer_8339 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_21063) ) ;
    buf_clk new_AGEMA_reg_buffer_8342 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T27), .Q (new_AGEMA_signal_21066) ) ;
    buf_clk new_AGEMA_reg_buffer_8345 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_21069) ) ;
    buf_clk new_AGEMA_reg_buffer_8348 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_21072) ) ;
    buf_clk new_AGEMA_reg_buffer_8351 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T10), .Q (new_AGEMA_signal_21075) ) ;
    buf_clk new_AGEMA_reg_buffer_8354 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_21078) ) ;
    buf_clk new_AGEMA_reg_buffer_8357 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_21081) ) ;
    buf_clk new_AGEMA_reg_buffer_8360 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T13), .Q (new_AGEMA_signal_21084) ) ;
    buf_clk new_AGEMA_reg_buffer_8363 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_21087) ) ;
    buf_clk new_AGEMA_reg_buffer_8366 ( .C (clk), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_21090) ) ;
    buf_clk new_AGEMA_reg_buffer_8369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T23), .Q (new_AGEMA_signal_21093) ) ;
    buf_clk new_AGEMA_reg_buffer_8372 ( .C (clk), .D (new_AGEMA_signal_6437), .Q (new_AGEMA_signal_21096) ) ;
    buf_clk new_AGEMA_reg_buffer_8375 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_21099) ) ;
    buf_clk new_AGEMA_reg_buffer_8378 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T19), .Q (new_AGEMA_signal_21102) ) ;
    buf_clk new_AGEMA_reg_buffer_8381 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_21105) ) ;
    buf_clk new_AGEMA_reg_buffer_8384 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_21108) ) ;
    buf_clk new_AGEMA_reg_buffer_8387 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T3), .Q (new_AGEMA_signal_21111) ) ;
    buf_clk new_AGEMA_reg_buffer_8390 ( .C (clk), .D (new_AGEMA_signal_5621), .Q (new_AGEMA_signal_21114) ) ;
    buf_clk new_AGEMA_reg_buffer_8393 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_21117) ) ;
    buf_clk new_AGEMA_reg_buffer_8396 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T22), .Q (new_AGEMA_signal_21120) ) ;
    buf_clk new_AGEMA_reg_buffer_8399 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_21123) ) ;
    buf_clk new_AGEMA_reg_buffer_8402 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_21126) ) ;
    buf_clk new_AGEMA_reg_buffer_8405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T20), .Q (new_AGEMA_signal_21129) ) ;
    buf_clk new_AGEMA_reg_buffer_8408 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_21132) ) ;
    buf_clk new_AGEMA_reg_buffer_8411 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_21135) ) ;
    buf_clk new_AGEMA_reg_buffer_8414 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T1), .Q (new_AGEMA_signal_21138) ) ;
    buf_clk new_AGEMA_reg_buffer_8417 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_21141) ) ;
    buf_clk new_AGEMA_reg_buffer_8420 ( .C (clk), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_21144) ) ;
    buf_clk new_AGEMA_reg_buffer_8423 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T4), .Q (new_AGEMA_signal_21147) ) ;
    buf_clk new_AGEMA_reg_buffer_8426 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_21150) ) ;
    buf_clk new_AGEMA_reg_buffer_8429 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_21153) ) ;
    buf_clk new_AGEMA_reg_buffer_8432 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_T2), .Q (new_AGEMA_signal_21156) ) ;
    buf_clk new_AGEMA_reg_buffer_8435 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_21159) ) ;
    buf_clk new_AGEMA_reg_buffer_8438 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_21162) ) ;
    buf_clk new_AGEMA_reg_buffer_8441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T6), .Q (new_AGEMA_signal_21165) ) ;
    buf_clk new_AGEMA_reg_buffer_8444 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_21168) ) ;
    buf_clk new_AGEMA_reg_buffer_8447 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_21171) ) ;
    buf_clk new_AGEMA_reg_buffer_8450 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T8), .Q (new_AGEMA_signal_21174) ) ;
    buf_clk new_AGEMA_reg_buffer_8453 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_21177) ) ;
    buf_clk new_AGEMA_reg_buffer_8456 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_21180) ) ;
    buf_clk new_AGEMA_reg_buffer_8459 ( .C (clk), .D (ciphertext_s0[96]), .Q (new_AGEMA_signal_21183) ) ;
    buf_clk new_AGEMA_reg_buffer_8462 ( .C (clk), .D (ciphertext_s1[96]), .Q (new_AGEMA_signal_21186) ) ;
    buf_clk new_AGEMA_reg_buffer_8465 ( .C (clk), .D (ciphertext_s2[96]), .Q (new_AGEMA_signal_21189) ) ;
    buf_clk new_AGEMA_reg_buffer_8468 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T16), .Q (new_AGEMA_signal_21192) ) ;
    buf_clk new_AGEMA_reg_buffer_8471 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_21195) ) ;
    buf_clk new_AGEMA_reg_buffer_8474 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_21198) ) ;
    buf_clk new_AGEMA_reg_buffer_8477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T9), .Q (new_AGEMA_signal_21201) ) ;
    buf_clk new_AGEMA_reg_buffer_8480 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_21204) ) ;
    buf_clk new_AGEMA_reg_buffer_8483 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_21207) ) ;
    buf_clk new_AGEMA_reg_buffer_8486 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T17), .Q (new_AGEMA_signal_21210) ) ;
    buf_clk new_AGEMA_reg_buffer_8489 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_21213) ) ;
    buf_clk new_AGEMA_reg_buffer_8492 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_21216) ) ;
    buf_clk new_AGEMA_reg_buffer_8495 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T15), .Q (new_AGEMA_signal_21219) ) ;
    buf_clk new_AGEMA_reg_buffer_8498 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_21222) ) ;
    buf_clk new_AGEMA_reg_buffer_8501 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_21225) ) ;
    buf_clk new_AGEMA_reg_buffer_8504 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T27), .Q (new_AGEMA_signal_21228) ) ;
    buf_clk new_AGEMA_reg_buffer_8507 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_21231) ) ;
    buf_clk new_AGEMA_reg_buffer_8510 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_21234) ) ;
    buf_clk new_AGEMA_reg_buffer_8513 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T10), .Q (new_AGEMA_signal_21237) ) ;
    buf_clk new_AGEMA_reg_buffer_8516 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_21240) ) ;
    buf_clk new_AGEMA_reg_buffer_8519 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_21243) ) ;
    buf_clk new_AGEMA_reg_buffer_8522 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T13), .Q (new_AGEMA_signal_21246) ) ;
    buf_clk new_AGEMA_reg_buffer_8525 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_21249) ) ;
    buf_clk new_AGEMA_reg_buffer_8528 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_21252) ) ;
    buf_clk new_AGEMA_reg_buffer_8531 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T23), .Q (new_AGEMA_signal_21255) ) ;
    buf_clk new_AGEMA_reg_buffer_8534 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_21258) ) ;
    buf_clk new_AGEMA_reg_buffer_8537 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_21261) ) ;
    buf_clk new_AGEMA_reg_buffer_8540 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T19), .Q (new_AGEMA_signal_21264) ) ;
    buf_clk new_AGEMA_reg_buffer_8543 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_21267) ) ;
    buf_clk new_AGEMA_reg_buffer_8546 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_21270) ) ;
    buf_clk new_AGEMA_reg_buffer_8549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T3), .Q (new_AGEMA_signal_21273) ) ;
    buf_clk new_AGEMA_reg_buffer_8552 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_21276) ) ;
    buf_clk new_AGEMA_reg_buffer_8555 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_21279) ) ;
    buf_clk new_AGEMA_reg_buffer_8558 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T22), .Q (new_AGEMA_signal_21282) ) ;
    buf_clk new_AGEMA_reg_buffer_8561 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_21285) ) ;
    buf_clk new_AGEMA_reg_buffer_8564 ( .C (clk), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_21288) ) ;
    buf_clk new_AGEMA_reg_buffer_8567 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T20), .Q (new_AGEMA_signal_21291) ) ;
    buf_clk new_AGEMA_reg_buffer_8570 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_21294) ) ;
    buf_clk new_AGEMA_reg_buffer_8573 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_21297) ) ;
    buf_clk new_AGEMA_reg_buffer_8576 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T1), .Q (new_AGEMA_signal_21300) ) ;
    buf_clk new_AGEMA_reg_buffer_8579 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_21303) ) ;
    buf_clk new_AGEMA_reg_buffer_8582 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_21306) ) ;
    buf_clk new_AGEMA_reg_buffer_8585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T4), .Q (new_AGEMA_signal_21309) ) ;
    buf_clk new_AGEMA_reg_buffer_8588 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_21312) ) ;
    buf_clk new_AGEMA_reg_buffer_8591 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_21315) ) ;
    buf_clk new_AGEMA_reg_buffer_8594 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_T2), .Q (new_AGEMA_signal_21318) ) ;
    buf_clk new_AGEMA_reg_buffer_8597 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_21321) ) ;
    buf_clk new_AGEMA_reg_buffer_8600 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_21324) ) ;
    buf_clk new_AGEMA_reg_buffer_8603 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T6), .Q (new_AGEMA_signal_21327) ) ;
    buf_clk new_AGEMA_reg_buffer_8606 ( .C (clk), .D (new_AGEMA_signal_5989), .Q (new_AGEMA_signal_21330) ) ;
    buf_clk new_AGEMA_reg_buffer_8609 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_21333) ) ;
    buf_clk new_AGEMA_reg_buffer_8612 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T8), .Q (new_AGEMA_signal_21336) ) ;
    buf_clk new_AGEMA_reg_buffer_8615 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_21339) ) ;
    buf_clk new_AGEMA_reg_buffer_8618 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_21342) ) ;
    buf_clk new_AGEMA_reg_buffer_8621 ( .C (clk), .D (ciphertext_s0[104]), .Q (new_AGEMA_signal_21345) ) ;
    buf_clk new_AGEMA_reg_buffer_8624 ( .C (clk), .D (ciphertext_s1[104]), .Q (new_AGEMA_signal_21348) ) ;
    buf_clk new_AGEMA_reg_buffer_8627 ( .C (clk), .D (ciphertext_s2[104]), .Q (new_AGEMA_signal_21351) ) ;
    buf_clk new_AGEMA_reg_buffer_8630 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T16), .Q (new_AGEMA_signal_21354) ) ;
    buf_clk new_AGEMA_reg_buffer_8633 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_21357) ) ;
    buf_clk new_AGEMA_reg_buffer_8636 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_21360) ) ;
    buf_clk new_AGEMA_reg_buffer_8639 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T9), .Q (new_AGEMA_signal_21363) ) ;
    buf_clk new_AGEMA_reg_buffer_8642 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_21366) ) ;
    buf_clk new_AGEMA_reg_buffer_8645 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_21369) ) ;
    buf_clk new_AGEMA_reg_buffer_8648 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T17), .Q (new_AGEMA_signal_21372) ) ;
    buf_clk new_AGEMA_reg_buffer_8651 ( .C (clk), .D (new_AGEMA_signal_6485), .Q (new_AGEMA_signal_21375) ) ;
    buf_clk new_AGEMA_reg_buffer_8654 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_21378) ) ;
    buf_clk new_AGEMA_reg_buffer_8657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T15), .Q (new_AGEMA_signal_21381) ) ;
    buf_clk new_AGEMA_reg_buffer_8660 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_21384) ) ;
    buf_clk new_AGEMA_reg_buffer_8663 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_21387) ) ;
    buf_clk new_AGEMA_reg_buffer_8666 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T27), .Q (new_AGEMA_signal_21390) ) ;
    buf_clk new_AGEMA_reg_buffer_8669 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_21393) ) ;
    buf_clk new_AGEMA_reg_buffer_8672 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_21396) ) ;
    buf_clk new_AGEMA_reg_buffer_8675 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T10), .Q (new_AGEMA_signal_21399) ) ;
    buf_clk new_AGEMA_reg_buffer_8678 ( .C (clk), .D (new_AGEMA_signal_6481), .Q (new_AGEMA_signal_21402) ) ;
    buf_clk new_AGEMA_reg_buffer_8681 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_21405) ) ;
    buf_clk new_AGEMA_reg_buffer_8684 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T13), .Q (new_AGEMA_signal_21408) ) ;
    buf_clk new_AGEMA_reg_buffer_8687 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_21411) ) ;
    buf_clk new_AGEMA_reg_buffer_8690 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_21414) ) ;
    buf_clk new_AGEMA_reg_buffer_8693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T23), .Q (new_AGEMA_signal_21417) ) ;
    buf_clk new_AGEMA_reg_buffer_8696 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_21420) ) ;
    buf_clk new_AGEMA_reg_buffer_8699 ( .C (clk), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_21423) ) ;
    buf_clk new_AGEMA_reg_buffer_8702 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T19), .Q (new_AGEMA_signal_21426) ) ;
    buf_clk new_AGEMA_reg_buffer_8705 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_21429) ) ;
    buf_clk new_AGEMA_reg_buffer_8708 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_21432) ) ;
    buf_clk new_AGEMA_reg_buffer_8711 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T3), .Q (new_AGEMA_signal_21435) ) ;
    buf_clk new_AGEMA_reg_buffer_8714 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_21438) ) ;
    buf_clk new_AGEMA_reg_buffer_8717 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_21441) ) ;
    buf_clk new_AGEMA_reg_buffer_8720 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T22), .Q (new_AGEMA_signal_21444) ) ;
    buf_clk new_AGEMA_reg_buffer_8723 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_21447) ) ;
    buf_clk new_AGEMA_reg_buffer_8726 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_21450) ) ;
    buf_clk new_AGEMA_reg_buffer_8729 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T20), .Q (new_AGEMA_signal_21453) ) ;
    buf_clk new_AGEMA_reg_buffer_8732 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_21456) ) ;
    buf_clk new_AGEMA_reg_buffer_8735 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_21459) ) ;
    buf_clk new_AGEMA_reg_buffer_8738 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T1), .Q (new_AGEMA_signal_21462) ) ;
    buf_clk new_AGEMA_reg_buffer_8741 ( .C (clk), .D (new_AGEMA_signal_5657), .Q (new_AGEMA_signal_21465) ) ;
    buf_clk new_AGEMA_reg_buffer_8744 ( .C (clk), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_21468) ) ;
    buf_clk new_AGEMA_reg_buffer_8747 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T4), .Q (new_AGEMA_signal_21471) ) ;
    buf_clk new_AGEMA_reg_buffer_8750 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_21474) ) ;
    buf_clk new_AGEMA_reg_buffer_8753 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_21477) ) ;
    buf_clk new_AGEMA_reg_buffer_8756 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_T2), .Q (new_AGEMA_signal_21480) ) ;
    buf_clk new_AGEMA_reg_buffer_8759 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_21483) ) ;
    buf_clk new_AGEMA_reg_buffer_8762 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_21486) ) ;
    buf_clk new_AGEMA_reg_buffer_8765 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T6), .Q (new_AGEMA_signal_21489) ) ;
    buf_clk new_AGEMA_reg_buffer_8768 ( .C (clk), .D (new_AGEMA_signal_6005), .Q (new_AGEMA_signal_21492) ) ;
    buf_clk new_AGEMA_reg_buffer_8771 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_21495) ) ;
    buf_clk new_AGEMA_reg_buffer_8774 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T8), .Q (new_AGEMA_signal_21498) ) ;
    buf_clk new_AGEMA_reg_buffer_8777 ( .C (clk), .D (new_AGEMA_signal_6505), .Q (new_AGEMA_signal_21501) ) ;
    buf_clk new_AGEMA_reg_buffer_8780 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_21504) ) ;
    buf_clk new_AGEMA_reg_buffer_8783 ( .C (clk), .D (ciphertext_s0[112]), .Q (new_AGEMA_signal_21507) ) ;
    buf_clk new_AGEMA_reg_buffer_8786 ( .C (clk), .D (ciphertext_s1[112]), .Q (new_AGEMA_signal_21510) ) ;
    buf_clk new_AGEMA_reg_buffer_8789 ( .C (clk), .D (ciphertext_s2[112]), .Q (new_AGEMA_signal_21513) ) ;
    buf_clk new_AGEMA_reg_buffer_8792 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T16), .Q (new_AGEMA_signal_21516) ) ;
    buf_clk new_AGEMA_reg_buffer_8795 ( .C (clk), .D (new_AGEMA_signal_6013), .Q (new_AGEMA_signal_21519) ) ;
    buf_clk new_AGEMA_reg_buffer_8798 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_21522) ) ;
    buf_clk new_AGEMA_reg_buffer_8801 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T9), .Q (new_AGEMA_signal_21525) ) ;
    buf_clk new_AGEMA_reg_buffer_8804 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_21528) ) ;
    buf_clk new_AGEMA_reg_buffer_8807 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_21531) ) ;
    buf_clk new_AGEMA_reg_buffer_8810 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T17), .Q (new_AGEMA_signal_21534) ) ;
    buf_clk new_AGEMA_reg_buffer_8813 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_21537) ) ;
    buf_clk new_AGEMA_reg_buffer_8816 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_21540) ) ;
    buf_clk new_AGEMA_reg_buffer_8819 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T15), .Q (new_AGEMA_signal_21543) ) ;
    buf_clk new_AGEMA_reg_buffer_8822 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_21546) ) ;
    buf_clk new_AGEMA_reg_buffer_8825 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_21549) ) ;
    buf_clk new_AGEMA_reg_buffer_8828 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T27), .Q (new_AGEMA_signal_21552) ) ;
    buf_clk new_AGEMA_reg_buffer_8831 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_21555) ) ;
    buf_clk new_AGEMA_reg_buffer_8834 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_21558) ) ;
    buf_clk new_AGEMA_reg_buffer_8837 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T10), .Q (new_AGEMA_signal_21561) ) ;
    buf_clk new_AGEMA_reg_buffer_8840 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_21564) ) ;
    buf_clk new_AGEMA_reg_buffer_8843 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_21567) ) ;
    buf_clk new_AGEMA_reg_buffer_8846 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T13), .Q (new_AGEMA_signal_21570) ) ;
    buf_clk new_AGEMA_reg_buffer_8849 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_21573) ) ;
    buf_clk new_AGEMA_reg_buffer_8852 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_21576) ) ;
    buf_clk new_AGEMA_reg_buffer_8855 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T23), .Q (new_AGEMA_signal_21579) ) ;
    buf_clk new_AGEMA_reg_buffer_8858 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_21582) ) ;
    buf_clk new_AGEMA_reg_buffer_8861 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_21585) ) ;
    buf_clk new_AGEMA_reg_buffer_8864 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T19), .Q (new_AGEMA_signal_21588) ) ;
    buf_clk new_AGEMA_reg_buffer_8867 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_21591) ) ;
    buf_clk new_AGEMA_reg_buffer_8870 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_21594) ) ;
    buf_clk new_AGEMA_reg_buffer_8873 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T3), .Q (new_AGEMA_signal_21597) ) ;
    buf_clk new_AGEMA_reg_buffer_8876 ( .C (clk), .D (new_AGEMA_signal_5681), .Q (new_AGEMA_signal_21600) ) ;
    buf_clk new_AGEMA_reg_buffer_8879 ( .C (clk), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_21603) ) ;
    buf_clk new_AGEMA_reg_buffer_8882 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T22), .Q (new_AGEMA_signal_21606) ) ;
    buf_clk new_AGEMA_reg_buffer_8885 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_21609) ) ;
    buf_clk new_AGEMA_reg_buffer_8888 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_21612) ) ;
    buf_clk new_AGEMA_reg_buffer_8891 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T20), .Q (new_AGEMA_signal_21615) ) ;
    buf_clk new_AGEMA_reg_buffer_8894 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_21618) ) ;
    buf_clk new_AGEMA_reg_buffer_8897 ( .C (clk), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_21621) ) ;
    buf_clk new_AGEMA_reg_buffer_8900 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T1), .Q (new_AGEMA_signal_21624) ) ;
    buf_clk new_AGEMA_reg_buffer_8903 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_21627) ) ;
    buf_clk new_AGEMA_reg_buffer_8906 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_21630) ) ;
    buf_clk new_AGEMA_reg_buffer_8909 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T4), .Q (new_AGEMA_signal_21633) ) ;
    buf_clk new_AGEMA_reg_buffer_8912 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_21636) ) ;
    buf_clk new_AGEMA_reg_buffer_8915 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_21639) ) ;
    buf_clk new_AGEMA_reg_buffer_8918 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_T2), .Q (new_AGEMA_signal_21642) ) ;
    buf_clk new_AGEMA_reg_buffer_8921 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_21645) ) ;
    buf_clk new_AGEMA_reg_buffer_8924 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_21648) ) ;
    buf_clk new_AGEMA_reg_buffer_8927 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T6), .Q (new_AGEMA_signal_21651) ) ;
    buf_clk new_AGEMA_reg_buffer_8930 ( .C (clk), .D (new_AGEMA_signal_6021), .Q (new_AGEMA_signal_21654) ) ;
    buf_clk new_AGEMA_reg_buffer_8933 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_21657) ) ;
    buf_clk new_AGEMA_reg_buffer_8936 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T8), .Q (new_AGEMA_signal_21660) ) ;
    buf_clk new_AGEMA_reg_buffer_8939 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_21663) ) ;
    buf_clk new_AGEMA_reg_buffer_8942 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_21666) ) ;
    buf_clk new_AGEMA_reg_buffer_8945 ( .C (clk), .D (ciphertext_s0[120]), .Q (new_AGEMA_signal_21669) ) ;
    buf_clk new_AGEMA_reg_buffer_8948 ( .C (clk), .D (ciphertext_s1[120]), .Q (new_AGEMA_signal_21672) ) ;
    buf_clk new_AGEMA_reg_buffer_8951 ( .C (clk), .D (ciphertext_s2[120]), .Q (new_AGEMA_signal_21675) ) ;
    buf_clk new_AGEMA_reg_buffer_8954 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T16), .Q (new_AGEMA_signal_21678) ) ;
    buf_clk new_AGEMA_reg_buffer_8957 ( .C (clk), .D (new_AGEMA_signal_6029), .Q (new_AGEMA_signal_21681) ) ;
    buf_clk new_AGEMA_reg_buffer_8960 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_21684) ) ;
    buf_clk new_AGEMA_reg_buffer_8963 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T9), .Q (new_AGEMA_signal_21687) ) ;
    buf_clk new_AGEMA_reg_buffer_8966 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_21690) ) ;
    buf_clk new_AGEMA_reg_buffer_8969 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_21693) ) ;
    buf_clk new_AGEMA_reg_buffer_8972 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T17), .Q (new_AGEMA_signal_21696) ) ;
    buf_clk new_AGEMA_reg_buffer_8975 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_21699) ) ;
    buf_clk new_AGEMA_reg_buffer_8978 ( .C (clk), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_21702) ) ;
    buf_clk new_AGEMA_reg_buffer_8981 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T15), .Q (new_AGEMA_signal_21705) ) ;
    buf_clk new_AGEMA_reg_buffer_8984 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_21708) ) ;
    buf_clk new_AGEMA_reg_buffer_8987 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_21711) ) ;
    buf_clk new_AGEMA_reg_buffer_8990 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T27), .Q (new_AGEMA_signal_21714) ) ;
    buf_clk new_AGEMA_reg_buffer_8993 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_21717) ) ;
    buf_clk new_AGEMA_reg_buffer_8996 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_21720) ) ;
    buf_clk new_AGEMA_reg_buffer_8999 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T10), .Q (new_AGEMA_signal_21723) ) ;
    buf_clk new_AGEMA_reg_buffer_9002 ( .C (clk), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_21726) ) ;
    buf_clk new_AGEMA_reg_buffer_9005 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_21729) ) ;
    buf_clk new_AGEMA_reg_buffer_9008 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T13), .Q (new_AGEMA_signal_21732) ) ;
    buf_clk new_AGEMA_reg_buffer_9011 ( .C (clk), .D (new_AGEMA_signal_6025), .Q (new_AGEMA_signal_21735) ) ;
    buf_clk new_AGEMA_reg_buffer_9014 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_21738) ) ;
    buf_clk new_AGEMA_reg_buffer_9017 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T23), .Q (new_AGEMA_signal_21741) ) ;
    buf_clk new_AGEMA_reg_buffer_9020 ( .C (clk), .D (new_AGEMA_signal_6541), .Q (new_AGEMA_signal_21744) ) ;
    buf_clk new_AGEMA_reg_buffer_9023 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_21747) ) ;
    buf_clk new_AGEMA_reg_buffer_9026 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T19), .Q (new_AGEMA_signal_21750) ) ;
    buf_clk new_AGEMA_reg_buffer_9029 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_21753) ) ;
    buf_clk new_AGEMA_reg_buffer_9032 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_21756) ) ;
    buf_clk new_AGEMA_reg_buffer_9035 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T3), .Q (new_AGEMA_signal_21759) ) ;
    buf_clk new_AGEMA_reg_buffer_9038 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_21762) ) ;
    buf_clk new_AGEMA_reg_buffer_9041 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_21765) ) ;
    buf_clk new_AGEMA_reg_buffer_9044 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T22), .Q (new_AGEMA_signal_21768) ) ;
    buf_clk new_AGEMA_reg_buffer_9047 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_21771) ) ;
    buf_clk new_AGEMA_reg_buffer_9050 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_21774) ) ;
    buf_clk new_AGEMA_reg_buffer_9053 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T20), .Q (new_AGEMA_signal_21777) ) ;
    buf_clk new_AGEMA_reg_buffer_9056 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_21780) ) ;
    buf_clk new_AGEMA_reg_buffer_9059 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_21783) ) ;
    buf_clk new_AGEMA_reg_buffer_9062 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T1), .Q (new_AGEMA_signal_21786) ) ;
    buf_clk new_AGEMA_reg_buffer_9065 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_21789) ) ;
    buf_clk new_AGEMA_reg_buffer_9068 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_21792) ) ;
    buf_clk new_AGEMA_reg_buffer_9071 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T4), .Q (new_AGEMA_signal_21795) ) ;
    buf_clk new_AGEMA_reg_buffer_9074 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_21798) ) ;
    buf_clk new_AGEMA_reg_buffer_9077 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_21801) ) ;
    buf_clk new_AGEMA_reg_buffer_9080 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_T2), .Q (new_AGEMA_signal_21804) ) ;
    buf_clk new_AGEMA_reg_buffer_9083 ( .C (clk), .D (new_AGEMA_signal_5699), .Q (new_AGEMA_signal_21807) ) ;
    buf_clk new_AGEMA_reg_buffer_9086 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_21810) ) ;
    buf_clk new_AGEMA_reg_buffer_9089 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_21813) ) ;
    buf_clk new_AGEMA_reg_buffer_9093 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_21817) ) ;
    buf_clk new_AGEMA_reg_buffer_9097 ( .C (clk), .D (key_s2[0]), .Q (new_AGEMA_signal_21821) ) ;
    buf_clk new_AGEMA_reg_buffer_9101 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_21825) ) ;
    buf_clk new_AGEMA_reg_buffer_9105 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_21829) ) ;
    buf_clk new_AGEMA_reg_buffer_9109 ( .C (clk), .D (key_s2[1]), .Q (new_AGEMA_signal_21833) ) ;
    buf_clk new_AGEMA_reg_buffer_9113 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_21837) ) ;
    buf_clk new_AGEMA_reg_buffer_9117 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_21841) ) ;
    buf_clk new_AGEMA_reg_buffer_9121 ( .C (clk), .D (key_s2[2]), .Q (new_AGEMA_signal_21845) ) ;
    buf_clk new_AGEMA_reg_buffer_9125 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_21849) ) ;
    buf_clk new_AGEMA_reg_buffer_9129 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_21853) ) ;
    buf_clk new_AGEMA_reg_buffer_9133 ( .C (clk), .D (key_s2[3]), .Q (new_AGEMA_signal_21857) ) ;
    buf_clk new_AGEMA_reg_buffer_9137 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_21861) ) ;
    buf_clk new_AGEMA_reg_buffer_9141 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_21865) ) ;
    buf_clk new_AGEMA_reg_buffer_9145 ( .C (clk), .D (key_s2[4]), .Q (new_AGEMA_signal_21869) ) ;
    buf_clk new_AGEMA_reg_buffer_9149 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_21873) ) ;
    buf_clk new_AGEMA_reg_buffer_9153 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_21877) ) ;
    buf_clk new_AGEMA_reg_buffer_9157 ( .C (clk), .D (key_s2[5]), .Q (new_AGEMA_signal_21881) ) ;
    buf_clk new_AGEMA_reg_buffer_9161 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_21885) ) ;
    buf_clk new_AGEMA_reg_buffer_9165 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_21889) ) ;
    buf_clk new_AGEMA_reg_buffer_9169 ( .C (clk), .D (key_s2[6]), .Q (new_AGEMA_signal_21893) ) ;
    buf_clk new_AGEMA_reg_buffer_9173 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_21897) ) ;
    buf_clk new_AGEMA_reg_buffer_9177 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_21901) ) ;
    buf_clk new_AGEMA_reg_buffer_9181 ( .C (clk), .D (key_s2[7]), .Q (new_AGEMA_signal_21905) ) ;
    buf_clk new_AGEMA_reg_buffer_9185 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_21909) ) ;
    buf_clk new_AGEMA_reg_buffer_9189 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_21913) ) ;
    buf_clk new_AGEMA_reg_buffer_9193 ( .C (clk), .D (key_s2[8]), .Q (new_AGEMA_signal_21917) ) ;
    buf_clk new_AGEMA_reg_buffer_9197 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_21921) ) ;
    buf_clk new_AGEMA_reg_buffer_9201 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_21925) ) ;
    buf_clk new_AGEMA_reg_buffer_9205 ( .C (clk), .D (key_s2[9]), .Q (new_AGEMA_signal_21929) ) ;
    buf_clk new_AGEMA_reg_buffer_9209 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_21933) ) ;
    buf_clk new_AGEMA_reg_buffer_9213 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_21937) ) ;
    buf_clk new_AGEMA_reg_buffer_9217 ( .C (clk), .D (key_s2[10]), .Q (new_AGEMA_signal_21941) ) ;
    buf_clk new_AGEMA_reg_buffer_9221 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_21945) ) ;
    buf_clk new_AGEMA_reg_buffer_9225 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_21949) ) ;
    buf_clk new_AGEMA_reg_buffer_9229 ( .C (clk), .D (key_s2[11]), .Q (new_AGEMA_signal_21953) ) ;
    buf_clk new_AGEMA_reg_buffer_9233 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_21957) ) ;
    buf_clk new_AGEMA_reg_buffer_9237 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_21961) ) ;
    buf_clk new_AGEMA_reg_buffer_9241 ( .C (clk), .D (key_s2[12]), .Q (new_AGEMA_signal_21965) ) ;
    buf_clk new_AGEMA_reg_buffer_9245 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_21969) ) ;
    buf_clk new_AGEMA_reg_buffer_9249 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_21973) ) ;
    buf_clk new_AGEMA_reg_buffer_9253 ( .C (clk), .D (key_s2[13]), .Q (new_AGEMA_signal_21977) ) ;
    buf_clk new_AGEMA_reg_buffer_9257 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_21981) ) ;
    buf_clk new_AGEMA_reg_buffer_9261 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_21985) ) ;
    buf_clk new_AGEMA_reg_buffer_9265 ( .C (clk), .D (key_s2[14]), .Q (new_AGEMA_signal_21989) ) ;
    buf_clk new_AGEMA_reg_buffer_9269 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_21993) ) ;
    buf_clk new_AGEMA_reg_buffer_9273 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_21997) ) ;
    buf_clk new_AGEMA_reg_buffer_9277 ( .C (clk), .D (key_s2[15]), .Q (new_AGEMA_signal_22001) ) ;
    buf_clk new_AGEMA_reg_buffer_9281 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_22005) ) ;
    buf_clk new_AGEMA_reg_buffer_9285 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_22009) ) ;
    buf_clk new_AGEMA_reg_buffer_9289 ( .C (clk), .D (key_s2[16]), .Q (new_AGEMA_signal_22013) ) ;
    buf_clk new_AGEMA_reg_buffer_9293 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_22017) ) ;
    buf_clk new_AGEMA_reg_buffer_9297 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_22021) ) ;
    buf_clk new_AGEMA_reg_buffer_9301 ( .C (clk), .D (key_s2[17]), .Q (new_AGEMA_signal_22025) ) ;
    buf_clk new_AGEMA_reg_buffer_9305 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_22029) ) ;
    buf_clk new_AGEMA_reg_buffer_9309 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_22033) ) ;
    buf_clk new_AGEMA_reg_buffer_9313 ( .C (clk), .D (key_s2[18]), .Q (new_AGEMA_signal_22037) ) ;
    buf_clk new_AGEMA_reg_buffer_9317 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_22041) ) ;
    buf_clk new_AGEMA_reg_buffer_9321 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_22045) ) ;
    buf_clk new_AGEMA_reg_buffer_9325 ( .C (clk), .D (key_s2[19]), .Q (new_AGEMA_signal_22049) ) ;
    buf_clk new_AGEMA_reg_buffer_9329 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_22053) ) ;
    buf_clk new_AGEMA_reg_buffer_9333 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_22057) ) ;
    buf_clk new_AGEMA_reg_buffer_9337 ( .C (clk), .D (key_s2[20]), .Q (new_AGEMA_signal_22061) ) ;
    buf_clk new_AGEMA_reg_buffer_9341 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_22065) ) ;
    buf_clk new_AGEMA_reg_buffer_9345 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_22069) ) ;
    buf_clk new_AGEMA_reg_buffer_9349 ( .C (clk), .D (key_s2[21]), .Q (new_AGEMA_signal_22073) ) ;
    buf_clk new_AGEMA_reg_buffer_9353 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_22077) ) ;
    buf_clk new_AGEMA_reg_buffer_9357 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_22081) ) ;
    buf_clk new_AGEMA_reg_buffer_9361 ( .C (clk), .D (key_s2[22]), .Q (new_AGEMA_signal_22085) ) ;
    buf_clk new_AGEMA_reg_buffer_9365 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_22089) ) ;
    buf_clk new_AGEMA_reg_buffer_9369 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_22093) ) ;
    buf_clk new_AGEMA_reg_buffer_9373 ( .C (clk), .D (key_s2[23]), .Q (new_AGEMA_signal_22097) ) ;
    buf_clk new_AGEMA_reg_buffer_9377 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_22101) ) ;
    buf_clk new_AGEMA_reg_buffer_9381 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_22105) ) ;
    buf_clk new_AGEMA_reg_buffer_9385 ( .C (clk), .D (key_s2[24]), .Q (new_AGEMA_signal_22109) ) ;
    buf_clk new_AGEMA_reg_buffer_9389 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_22113) ) ;
    buf_clk new_AGEMA_reg_buffer_9393 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_22117) ) ;
    buf_clk new_AGEMA_reg_buffer_9397 ( .C (clk), .D (key_s2[25]), .Q (new_AGEMA_signal_22121) ) ;
    buf_clk new_AGEMA_reg_buffer_9401 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_22125) ) ;
    buf_clk new_AGEMA_reg_buffer_9405 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_22129) ) ;
    buf_clk new_AGEMA_reg_buffer_9409 ( .C (clk), .D (key_s2[26]), .Q (new_AGEMA_signal_22133) ) ;
    buf_clk new_AGEMA_reg_buffer_9413 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_22137) ) ;
    buf_clk new_AGEMA_reg_buffer_9417 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_22141) ) ;
    buf_clk new_AGEMA_reg_buffer_9421 ( .C (clk), .D (key_s2[27]), .Q (new_AGEMA_signal_22145) ) ;
    buf_clk new_AGEMA_reg_buffer_9425 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_22149) ) ;
    buf_clk new_AGEMA_reg_buffer_9429 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_22153) ) ;
    buf_clk new_AGEMA_reg_buffer_9433 ( .C (clk), .D (key_s2[28]), .Q (new_AGEMA_signal_22157) ) ;
    buf_clk new_AGEMA_reg_buffer_9437 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_22161) ) ;
    buf_clk new_AGEMA_reg_buffer_9441 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_22165) ) ;
    buf_clk new_AGEMA_reg_buffer_9445 ( .C (clk), .D (key_s2[29]), .Q (new_AGEMA_signal_22169) ) ;
    buf_clk new_AGEMA_reg_buffer_9449 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_22173) ) ;
    buf_clk new_AGEMA_reg_buffer_9453 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_22177) ) ;
    buf_clk new_AGEMA_reg_buffer_9457 ( .C (clk), .D (key_s2[30]), .Q (new_AGEMA_signal_22181) ) ;
    buf_clk new_AGEMA_reg_buffer_9461 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_22185) ) ;
    buf_clk new_AGEMA_reg_buffer_9465 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_22189) ) ;
    buf_clk new_AGEMA_reg_buffer_9469 ( .C (clk), .D (key_s2[31]), .Q (new_AGEMA_signal_22193) ) ;
    buf_clk new_AGEMA_reg_buffer_9473 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_22197) ) ;
    buf_clk new_AGEMA_reg_buffer_9477 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_22201) ) ;
    buf_clk new_AGEMA_reg_buffer_9481 ( .C (clk), .D (key_s2[32]), .Q (new_AGEMA_signal_22205) ) ;
    buf_clk new_AGEMA_reg_buffer_9485 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_22209) ) ;
    buf_clk new_AGEMA_reg_buffer_9489 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_22213) ) ;
    buf_clk new_AGEMA_reg_buffer_9493 ( .C (clk), .D (key_s2[33]), .Q (new_AGEMA_signal_22217) ) ;
    buf_clk new_AGEMA_reg_buffer_9497 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_22221) ) ;
    buf_clk new_AGEMA_reg_buffer_9501 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_22225) ) ;
    buf_clk new_AGEMA_reg_buffer_9505 ( .C (clk), .D (key_s2[34]), .Q (new_AGEMA_signal_22229) ) ;
    buf_clk new_AGEMA_reg_buffer_9509 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_22233) ) ;
    buf_clk new_AGEMA_reg_buffer_9513 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_22237) ) ;
    buf_clk new_AGEMA_reg_buffer_9517 ( .C (clk), .D (key_s2[35]), .Q (new_AGEMA_signal_22241) ) ;
    buf_clk new_AGEMA_reg_buffer_9521 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_22245) ) ;
    buf_clk new_AGEMA_reg_buffer_9525 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_22249) ) ;
    buf_clk new_AGEMA_reg_buffer_9529 ( .C (clk), .D (key_s2[36]), .Q (new_AGEMA_signal_22253) ) ;
    buf_clk new_AGEMA_reg_buffer_9533 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_22257) ) ;
    buf_clk new_AGEMA_reg_buffer_9537 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_22261) ) ;
    buf_clk new_AGEMA_reg_buffer_9541 ( .C (clk), .D (key_s2[37]), .Q (new_AGEMA_signal_22265) ) ;
    buf_clk new_AGEMA_reg_buffer_9545 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_22269) ) ;
    buf_clk new_AGEMA_reg_buffer_9549 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_22273) ) ;
    buf_clk new_AGEMA_reg_buffer_9553 ( .C (clk), .D (key_s2[38]), .Q (new_AGEMA_signal_22277) ) ;
    buf_clk new_AGEMA_reg_buffer_9557 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_22281) ) ;
    buf_clk new_AGEMA_reg_buffer_9561 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_22285) ) ;
    buf_clk new_AGEMA_reg_buffer_9565 ( .C (clk), .D (key_s2[39]), .Q (new_AGEMA_signal_22289) ) ;
    buf_clk new_AGEMA_reg_buffer_9569 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_22293) ) ;
    buf_clk new_AGEMA_reg_buffer_9573 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_22297) ) ;
    buf_clk new_AGEMA_reg_buffer_9577 ( .C (clk), .D (key_s2[40]), .Q (new_AGEMA_signal_22301) ) ;
    buf_clk new_AGEMA_reg_buffer_9581 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_22305) ) ;
    buf_clk new_AGEMA_reg_buffer_9585 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_22309) ) ;
    buf_clk new_AGEMA_reg_buffer_9589 ( .C (clk), .D (key_s2[41]), .Q (new_AGEMA_signal_22313) ) ;
    buf_clk new_AGEMA_reg_buffer_9593 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_22317) ) ;
    buf_clk new_AGEMA_reg_buffer_9597 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_22321) ) ;
    buf_clk new_AGEMA_reg_buffer_9601 ( .C (clk), .D (key_s2[42]), .Q (new_AGEMA_signal_22325) ) ;
    buf_clk new_AGEMA_reg_buffer_9605 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_22329) ) ;
    buf_clk new_AGEMA_reg_buffer_9609 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_22333) ) ;
    buf_clk new_AGEMA_reg_buffer_9613 ( .C (clk), .D (key_s2[43]), .Q (new_AGEMA_signal_22337) ) ;
    buf_clk new_AGEMA_reg_buffer_9617 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_22341) ) ;
    buf_clk new_AGEMA_reg_buffer_9621 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_22345) ) ;
    buf_clk new_AGEMA_reg_buffer_9625 ( .C (clk), .D (key_s2[44]), .Q (new_AGEMA_signal_22349) ) ;
    buf_clk new_AGEMA_reg_buffer_9629 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_22353) ) ;
    buf_clk new_AGEMA_reg_buffer_9633 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_22357) ) ;
    buf_clk new_AGEMA_reg_buffer_9637 ( .C (clk), .D (key_s2[45]), .Q (new_AGEMA_signal_22361) ) ;
    buf_clk new_AGEMA_reg_buffer_9641 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_22365) ) ;
    buf_clk new_AGEMA_reg_buffer_9645 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_22369) ) ;
    buf_clk new_AGEMA_reg_buffer_9649 ( .C (clk), .D (key_s2[46]), .Q (new_AGEMA_signal_22373) ) ;
    buf_clk new_AGEMA_reg_buffer_9653 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_22377) ) ;
    buf_clk new_AGEMA_reg_buffer_9657 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_22381) ) ;
    buf_clk new_AGEMA_reg_buffer_9661 ( .C (clk), .D (key_s2[47]), .Q (new_AGEMA_signal_22385) ) ;
    buf_clk new_AGEMA_reg_buffer_9665 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_22389) ) ;
    buf_clk new_AGEMA_reg_buffer_9669 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_22393) ) ;
    buf_clk new_AGEMA_reg_buffer_9673 ( .C (clk), .D (key_s2[48]), .Q (new_AGEMA_signal_22397) ) ;
    buf_clk new_AGEMA_reg_buffer_9677 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_22401) ) ;
    buf_clk new_AGEMA_reg_buffer_9681 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_22405) ) ;
    buf_clk new_AGEMA_reg_buffer_9685 ( .C (clk), .D (key_s2[49]), .Q (new_AGEMA_signal_22409) ) ;
    buf_clk new_AGEMA_reg_buffer_9689 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_22413) ) ;
    buf_clk new_AGEMA_reg_buffer_9693 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_22417) ) ;
    buf_clk new_AGEMA_reg_buffer_9697 ( .C (clk), .D (key_s2[50]), .Q (new_AGEMA_signal_22421) ) ;
    buf_clk new_AGEMA_reg_buffer_9701 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_22425) ) ;
    buf_clk new_AGEMA_reg_buffer_9705 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_22429) ) ;
    buf_clk new_AGEMA_reg_buffer_9709 ( .C (clk), .D (key_s2[51]), .Q (new_AGEMA_signal_22433) ) ;
    buf_clk new_AGEMA_reg_buffer_9713 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_22437) ) ;
    buf_clk new_AGEMA_reg_buffer_9717 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_22441) ) ;
    buf_clk new_AGEMA_reg_buffer_9721 ( .C (clk), .D (key_s2[52]), .Q (new_AGEMA_signal_22445) ) ;
    buf_clk new_AGEMA_reg_buffer_9725 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_22449) ) ;
    buf_clk new_AGEMA_reg_buffer_9729 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_22453) ) ;
    buf_clk new_AGEMA_reg_buffer_9733 ( .C (clk), .D (key_s2[53]), .Q (new_AGEMA_signal_22457) ) ;
    buf_clk new_AGEMA_reg_buffer_9737 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_22461) ) ;
    buf_clk new_AGEMA_reg_buffer_9741 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_22465) ) ;
    buf_clk new_AGEMA_reg_buffer_9745 ( .C (clk), .D (key_s2[54]), .Q (new_AGEMA_signal_22469) ) ;
    buf_clk new_AGEMA_reg_buffer_9749 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_22473) ) ;
    buf_clk new_AGEMA_reg_buffer_9753 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_22477) ) ;
    buf_clk new_AGEMA_reg_buffer_9757 ( .C (clk), .D (key_s2[55]), .Q (new_AGEMA_signal_22481) ) ;
    buf_clk new_AGEMA_reg_buffer_9761 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_22485) ) ;
    buf_clk new_AGEMA_reg_buffer_9765 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_22489) ) ;
    buf_clk new_AGEMA_reg_buffer_9769 ( .C (clk), .D (key_s2[56]), .Q (new_AGEMA_signal_22493) ) ;
    buf_clk new_AGEMA_reg_buffer_9773 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_22497) ) ;
    buf_clk new_AGEMA_reg_buffer_9777 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_22501) ) ;
    buf_clk new_AGEMA_reg_buffer_9781 ( .C (clk), .D (key_s2[57]), .Q (new_AGEMA_signal_22505) ) ;
    buf_clk new_AGEMA_reg_buffer_9785 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_22509) ) ;
    buf_clk new_AGEMA_reg_buffer_9789 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_22513) ) ;
    buf_clk new_AGEMA_reg_buffer_9793 ( .C (clk), .D (key_s2[58]), .Q (new_AGEMA_signal_22517) ) ;
    buf_clk new_AGEMA_reg_buffer_9797 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_22521) ) ;
    buf_clk new_AGEMA_reg_buffer_9801 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_22525) ) ;
    buf_clk new_AGEMA_reg_buffer_9805 ( .C (clk), .D (key_s2[59]), .Q (new_AGEMA_signal_22529) ) ;
    buf_clk new_AGEMA_reg_buffer_9809 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_22533) ) ;
    buf_clk new_AGEMA_reg_buffer_9813 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_22537) ) ;
    buf_clk new_AGEMA_reg_buffer_9817 ( .C (clk), .D (key_s2[60]), .Q (new_AGEMA_signal_22541) ) ;
    buf_clk new_AGEMA_reg_buffer_9821 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_22545) ) ;
    buf_clk new_AGEMA_reg_buffer_9825 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_22549) ) ;
    buf_clk new_AGEMA_reg_buffer_9829 ( .C (clk), .D (key_s2[61]), .Q (new_AGEMA_signal_22553) ) ;
    buf_clk new_AGEMA_reg_buffer_9833 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_22557) ) ;
    buf_clk new_AGEMA_reg_buffer_9837 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_22561) ) ;
    buf_clk new_AGEMA_reg_buffer_9841 ( .C (clk), .D (key_s2[62]), .Q (new_AGEMA_signal_22565) ) ;
    buf_clk new_AGEMA_reg_buffer_9845 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_22569) ) ;
    buf_clk new_AGEMA_reg_buffer_9849 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_22573) ) ;
    buf_clk new_AGEMA_reg_buffer_9853 ( .C (clk), .D (key_s2[63]), .Q (new_AGEMA_signal_22577) ) ;
    buf_clk new_AGEMA_reg_buffer_9857 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_22581) ) ;
    buf_clk new_AGEMA_reg_buffer_9861 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_22585) ) ;
    buf_clk new_AGEMA_reg_buffer_9865 ( .C (clk), .D (key_s2[64]), .Q (new_AGEMA_signal_22589) ) ;
    buf_clk new_AGEMA_reg_buffer_9869 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_22593) ) ;
    buf_clk new_AGEMA_reg_buffer_9873 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_22597) ) ;
    buf_clk new_AGEMA_reg_buffer_9877 ( .C (clk), .D (key_s2[65]), .Q (new_AGEMA_signal_22601) ) ;
    buf_clk new_AGEMA_reg_buffer_9881 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_22605) ) ;
    buf_clk new_AGEMA_reg_buffer_9885 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_22609) ) ;
    buf_clk new_AGEMA_reg_buffer_9889 ( .C (clk), .D (key_s2[66]), .Q (new_AGEMA_signal_22613) ) ;
    buf_clk new_AGEMA_reg_buffer_9893 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_22617) ) ;
    buf_clk new_AGEMA_reg_buffer_9897 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_22621) ) ;
    buf_clk new_AGEMA_reg_buffer_9901 ( .C (clk), .D (key_s2[67]), .Q (new_AGEMA_signal_22625) ) ;
    buf_clk new_AGEMA_reg_buffer_9905 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_22629) ) ;
    buf_clk new_AGEMA_reg_buffer_9909 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_22633) ) ;
    buf_clk new_AGEMA_reg_buffer_9913 ( .C (clk), .D (key_s2[68]), .Q (new_AGEMA_signal_22637) ) ;
    buf_clk new_AGEMA_reg_buffer_9917 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_22641) ) ;
    buf_clk new_AGEMA_reg_buffer_9921 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_22645) ) ;
    buf_clk new_AGEMA_reg_buffer_9925 ( .C (clk), .D (key_s2[69]), .Q (new_AGEMA_signal_22649) ) ;
    buf_clk new_AGEMA_reg_buffer_9929 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_22653) ) ;
    buf_clk new_AGEMA_reg_buffer_9933 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_22657) ) ;
    buf_clk new_AGEMA_reg_buffer_9937 ( .C (clk), .D (key_s2[70]), .Q (new_AGEMA_signal_22661) ) ;
    buf_clk new_AGEMA_reg_buffer_9941 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_22665) ) ;
    buf_clk new_AGEMA_reg_buffer_9945 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_22669) ) ;
    buf_clk new_AGEMA_reg_buffer_9949 ( .C (clk), .D (key_s2[71]), .Q (new_AGEMA_signal_22673) ) ;
    buf_clk new_AGEMA_reg_buffer_9953 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_22677) ) ;
    buf_clk new_AGEMA_reg_buffer_9957 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_22681) ) ;
    buf_clk new_AGEMA_reg_buffer_9961 ( .C (clk), .D (key_s2[72]), .Q (new_AGEMA_signal_22685) ) ;
    buf_clk new_AGEMA_reg_buffer_9965 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_22689) ) ;
    buf_clk new_AGEMA_reg_buffer_9969 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_22693) ) ;
    buf_clk new_AGEMA_reg_buffer_9973 ( .C (clk), .D (key_s2[73]), .Q (new_AGEMA_signal_22697) ) ;
    buf_clk new_AGEMA_reg_buffer_9977 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_22701) ) ;
    buf_clk new_AGEMA_reg_buffer_9981 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_22705) ) ;
    buf_clk new_AGEMA_reg_buffer_9985 ( .C (clk), .D (key_s2[74]), .Q (new_AGEMA_signal_22709) ) ;
    buf_clk new_AGEMA_reg_buffer_9989 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_22713) ) ;
    buf_clk new_AGEMA_reg_buffer_9993 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_22717) ) ;
    buf_clk new_AGEMA_reg_buffer_9997 ( .C (clk), .D (key_s2[75]), .Q (new_AGEMA_signal_22721) ) ;
    buf_clk new_AGEMA_reg_buffer_10001 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_22725) ) ;
    buf_clk new_AGEMA_reg_buffer_10005 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_22729) ) ;
    buf_clk new_AGEMA_reg_buffer_10009 ( .C (clk), .D (key_s2[76]), .Q (new_AGEMA_signal_22733) ) ;
    buf_clk new_AGEMA_reg_buffer_10013 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_22737) ) ;
    buf_clk new_AGEMA_reg_buffer_10017 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_22741) ) ;
    buf_clk new_AGEMA_reg_buffer_10021 ( .C (clk), .D (key_s2[77]), .Q (new_AGEMA_signal_22745) ) ;
    buf_clk new_AGEMA_reg_buffer_10025 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_22749) ) ;
    buf_clk new_AGEMA_reg_buffer_10029 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_22753) ) ;
    buf_clk new_AGEMA_reg_buffer_10033 ( .C (clk), .D (key_s2[78]), .Q (new_AGEMA_signal_22757) ) ;
    buf_clk new_AGEMA_reg_buffer_10037 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_22761) ) ;
    buf_clk new_AGEMA_reg_buffer_10041 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_22765) ) ;
    buf_clk new_AGEMA_reg_buffer_10045 ( .C (clk), .D (key_s2[79]), .Q (new_AGEMA_signal_22769) ) ;
    buf_clk new_AGEMA_reg_buffer_10049 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_22773) ) ;
    buf_clk new_AGEMA_reg_buffer_10053 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_22777) ) ;
    buf_clk new_AGEMA_reg_buffer_10057 ( .C (clk), .D (key_s2[80]), .Q (new_AGEMA_signal_22781) ) ;
    buf_clk new_AGEMA_reg_buffer_10061 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_22785) ) ;
    buf_clk new_AGEMA_reg_buffer_10065 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_22789) ) ;
    buf_clk new_AGEMA_reg_buffer_10069 ( .C (clk), .D (key_s2[81]), .Q (new_AGEMA_signal_22793) ) ;
    buf_clk new_AGEMA_reg_buffer_10073 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_22797) ) ;
    buf_clk new_AGEMA_reg_buffer_10077 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_22801) ) ;
    buf_clk new_AGEMA_reg_buffer_10081 ( .C (clk), .D (key_s2[82]), .Q (new_AGEMA_signal_22805) ) ;
    buf_clk new_AGEMA_reg_buffer_10085 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_22809) ) ;
    buf_clk new_AGEMA_reg_buffer_10089 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_22813) ) ;
    buf_clk new_AGEMA_reg_buffer_10093 ( .C (clk), .D (key_s2[83]), .Q (new_AGEMA_signal_22817) ) ;
    buf_clk new_AGEMA_reg_buffer_10097 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_22821) ) ;
    buf_clk new_AGEMA_reg_buffer_10101 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_22825) ) ;
    buf_clk new_AGEMA_reg_buffer_10105 ( .C (clk), .D (key_s2[84]), .Q (new_AGEMA_signal_22829) ) ;
    buf_clk new_AGEMA_reg_buffer_10109 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_22833) ) ;
    buf_clk new_AGEMA_reg_buffer_10113 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_22837) ) ;
    buf_clk new_AGEMA_reg_buffer_10117 ( .C (clk), .D (key_s2[85]), .Q (new_AGEMA_signal_22841) ) ;
    buf_clk new_AGEMA_reg_buffer_10121 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_22845) ) ;
    buf_clk new_AGEMA_reg_buffer_10125 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_22849) ) ;
    buf_clk new_AGEMA_reg_buffer_10129 ( .C (clk), .D (key_s2[86]), .Q (new_AGEMA_signal_22853) ) ;
    buf_clk new_AGEMA_reg_buffer_10133 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_22857) ) ;
    buf_clk new_AGEMA_reg_buffer_10137 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_22861) ) ;
    buf_clk new_AGEMA_reg_buffer_10141 ( .C (clk), .D (key_s2[87]), .Q (new_AGEMA_signal_22865) ) ;
    buf_clk new_AGEMA_reg_buffer_10145 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_22869) ) ;
    buf_clk new_AGEMA_reg_buffer_10149 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_22873) ) ;
    buf_clk new_AGEMA_reg_buffer_10153 ( .C (clk), .D (key_s2[88]), .Q (new_AGEMA_signal_22877) ) ;
    buf_clk new_AGEMA_reg_buffer_10157 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_22881) ) ;
    buf_clk new_AGEMA_reg_buffer_10161 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_22885) ) ;
    buf_clk new_AGEMA_reg_buffer_10165 ( .C (clk), .D (key_s2[89]), .Q (new_AGEMA_signal_22889) ) ;
    buf_clk new_AGEMA_reg_buffer_10169 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_22893) ) ;
    buf_clk new_AGEMA_reg_buffer_10173 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_22897) ) ;
    buf_clk new_AGEMA_reg_buffer_10177 ( .C (clk), .D (key_s2[90]), .Q (new_AGEMA_signal_22901) ) ;
    buf_clk new_AGEMA_reg_buffer_10181 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_22905) ) ;
    buf_clk new_AGEMA_reg_buffer_10185 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_22909) ) ;
    buf_clk new_AGEMA_reg_buffer_10189 ( .C (clk), .D (key_s2[91]), .Q (new_AGEMA_signal_22913) ) ;
    buf_clk new_AGEMA_reg_buffer_10193 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_22917) ) ;
    buf_clk new_AGEMA_reg_buffer_10197 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_22921) ) ;
    buf_clk new_AGEMA_reg_buffer_10201 ( .C (clk), .D (key_s2[92]), .Q (new_AGEMA_signal_22925) ) ;
    buf_clk new_AGEMA_reg_buffer_10205 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_22929) ) ;
    buf_clk new_AGEMA_reg_buffer_10209 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_22933) ) ;
    buf_clk new_AGEMA_reg_buffer_10213 ( .C (clk), .D (key_s2[93]), .Q (new_AGEMA_signal_22937) ) ;
    buf_clk new_AGEMA_reg_buffer_10217 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_22941) ) ;
    buf_clk new_AGEMA_reg_buffer_10221 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_22945) ) ;
    buf_clk new_AGEMA_reg_buffer_10225 ( .C (clk), .D (key_s2[94]), .Q (new_AGEMA_signal_22949) ) ;
    buf_clk new_AGEMA_reg_buffer_10229 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_22953) ) ;
    buf_clk new_AGEMA_reg_buffer_10233 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_22957) ) ;
    buf_clk new_AGEMA_reg_buffer_10237 ( .C (clk), .D (key_s2[95]), .Q (new_AGEMA_signal_22961) ) ;
    buf_clk new_AGEMA_reg_buffer_10241 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_22965) ) ;
    buf_clk new_AGEMA_reg_buffer_10245 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_22969) ) ;
    buf_clk new_AGEMA_reg_buffer_10249 ( .C (clk), .D (key_s2[96]), .Q (new_AGEMA_signal_22973) ) ;
    buf_clk new_AGEMA_reg_buffer_10253 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_22977) ) ;
    buf_clk new_AGEMA_reg_buffer_10257 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_22981) ) ;
    buf_clk new_AGEMA_reg_buffer_10261 ( .C (clk), .D (key_s2[97]), .Q (new_AGEMA_signal_22985) ) ;
    buf_clk new_AGEMA_reg_buffer_10265 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_22989) ) ;
    buf_clk new_AGEMA_reg_buffer_10269 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_22993) ) ;
    buf_clk new_AGEMA_reg_buffer_10273 ( .C (clk), .D (key_s2[98]), .Q (new_AGEMA_signal_22997) ) ;
    buf_clk new_AGEMA_reg_buffer_10277 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_23001) ) ;
    buf_clk new_AGEMA_reg_buffer_10281 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_23005) ) ;
    buf_clk new_AGEMA_reg_buffer_10285 ( .C (clk), .D (key_s2[99]), .Q (new_AGEMA_signal_23009) ) ;
    buf_clk new_AGEMA_reg_buffer_10289 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_23013) ) ;
    buf_clk new_AGEMA_reg_buffer_10293 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_23017) ) ;
    buf_clk new_AGEMA_reg_buffer_10297 ( .C (clk), .D (key_s2[100]), .Q (new_AGEMA_signal_23021) ) ;
    buf_clk new_AGEMA_reg_buffer_10301 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_23025) ) ;
    buf_clk new_AGEMA_reg_buffer_10305 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_23029) ) ;
    buf_clk new_AGEMA_reg_buffer_10309 ( .C (clk), .D (key_s2[101]), .Q (new_AGEMA_signal_23033) ) ;
    buf_clk new_AGEMA_reg_buffer_10313 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_23037) ) ;
    buf_clk new_AGEMA_reg_buffer_10317 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_23041) ) ;
    buf_clk new_AGEMA_reg_buffer_10321 ( .C (clk), .D (key_s2[102]), .Q (new_AGEMA_signal_23045) ) ;
    buf_clk new_AGEMA_reg_buffer_10325 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_23049) ) ;
    buf_clk new_AGEMA_reg_buffer_10329 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_23053) ) ;
    buf_clk new_AGEMA_reg_buffer_10333 ( .C (clk), .D (key_s2[103]), .Q (new_AGEMA_signal_23057) ) ;
    buf_clk new_AGEMA_reg_buffer_10337 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_23061) ) ;
    buf_clk new_AGEMA_reg_buffer_10341 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_23065) ) ;
    buf_clk new_AGEMA_reg_buffer_10345 ( .C (clk), .D (key_s2[104]), .Q (new_AGEMA_signal_23069) ) ;
    buf_clk new_AGEMA_reg_buffer_10349 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_23073) ) ;
    buf_clk new_AGEMA_reg_buffer_10353 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_23077) ) ;
    buf_clk new_AGEMA_reg_buffer_10357 ( .C (clk), .D (key_s2[105]), .Q (new_AGEMA_signal_23081) ) ;
    buf_clk new_AGEMA_reg_buffer_10361 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_23085) ) ;
    buf_clk new_AGEMA_reg_buffer_10365 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_23089) ) ;
    buf_clk new_AGEMA_reg_buffer_10369 ( .C (clk), .D (key_s2[106]), .Q (new_AGEMA_signal_23093) ) ;
    buf_clk new_AGEMA_reg_buffer_10373 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_23097) ) ;
    buf_clk new_AGEMA_reg_buffer_10377 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_23101) ) ;
    buf_clk new_AGEMA_reg_buffer_10381 ( .C (clk), .D (key_s2[107]), .Q (new_AGEMA_signal_23105) ) ;
    buf_clk new_AGEMA_reg_buffer_10385 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_23109) ) ;
    buf_clk new_AGEMA_reg_buffer_10389 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_23113) ) ;
    buf_clk new_AGEMA_reg_buffer_10393 ( .C (clk), .D (key_s2[108]), .Q (new_AGEMA_signal_23117) ) ;
    buf_clk new_AGEMA_reg_buffer_10397 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_23121) ) ;
    buf_clk new_AGEMA_reg_buffer_10401 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_23125) ) ;
    buf_clk new_AGEMA_reg_buffer_10405 ( .C (clk), .D (key_s2[109]), .Q (new_AGEMA_signal_23129) ) ;
    buf_clk new_AGEMA_reg_buffer_10409 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_23133) ) ;
    buf_clk new_AGEMA_reg_buffer_10413 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_23137) ) ;
    buf_clk new_AGEMA_reg_buffer_10417 ( .C (clk), .D (key_s2[110]), .Q (new_AGEMA_signal_23141) ) ;
    buf_clk new_AGEMA_reg_buffer_10421 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_23145) ) ;
    buf_clk new_AGEMA_reg_buffer_10425 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_23149) ) ;
    buf_clk new_AGEMA_reg_buffer_10429 ( .C (clk), .D (key_s2[111]), .Q (new_AGEMA_signal_23153) ) ;
    buf_clk new_AGEMA_reg_buffer_10433 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_23157) ) ;
    buf_clk new_AGEMA_reg_buffer_10437 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_23161) ) ;
    buf_clk new_AGEMA_reg_buffer_10441 ( .C (clk), .D (key_s2[112]), .Q (new_AGEMA_signal_23165) ) ;
    buf_clk new_AGEMA_reg_buffer_10445 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_23169) ) ;
    buf_clk new_AGEMA_reg_buffer_10449 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_23173) ) ;
    buf_clk new_AGEMA_reg_buffer_10453 ( .C (clk), .D (key_s2[113]), .Q (new_AGEMA_signal_23177) ) ;
    buf_clk new_AGEMA_reg_buffer_10457 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_23181) ) ;
    buf_clk new_AGEMA_reg_buffer_10461 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_23185) ) ;
    buf_clk new_AGEMA_reg_buffer_10465 ( .C (clk), .D (key_s2[114]), .Q (new_AGEMA_signal_23189) ) ;
    buf_clk new_AGEMA_reg_buffer_10469 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_23193) ) ;
    buf_clk new_AGEMA_reg_buffer_10473 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_23197) ) ;
    buf_clk new_AGEMA_reg_buffer_10477 ( .C (clk), .D (key_s2[115]), .Q (new_AGEMA_signal_23201) ) ;
    buf_clk new_AGEMA_reg_buffer_10481 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_23205) ) ;
    buf_clk new_AGEMA_reg_buffer_10485 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_23209) ) ;
    buf_clk new_AGEMA_reg_buffer_10489 ( .C (clk), .D (key_s2[116]), .Q (new_AGEMA_signal_23213) ) ;
    buf_clk new_AGEMA_reg_buffer_10493 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_23217) ) ;
    buf_clk new_AGEMA_reg_buffer_10497 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_23221) ) ;
    buf_clk new_AGEMA_reg_buffer_10501 ( .C (clk), .D (key_s2[117]), .Q (new_AGEMA_signal_23225) ) ;
    buf_clk new_AGEMA_reg_buffer_10505 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_23229) ) ;
    buf_clk new_AGEMA_reg_buffer_10509 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_23233) ) ;
    buf_clk new_AGEMA_reg_buffer_10513 ( .C (clk), .D (key_s2[118]), .Q (new_AGEMA_signal_23237) ) ;
    buf_clk new_AGEMA_reg_buffer_10517 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_23241) ) ;
    buf_clk new_AGEMA_reg_buffer_10521 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_23245) ) ;
    buf_clk new_AGEMA_reg_buffer_10525 ( .C (clk), .D (key_s2[119]), .Q (new_AGEMA_signal_23249) ) ;
    buf_clk new_AGEMA_reg_buffer_10529 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_23253) ) ;
    buf_clk new_AGEMA_reg_buffer_10533 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_23257) ) ;
    buf_clk new_AGEMA_reg_buffer_10537 ( .C (clk), .D (key_s2[120]), .Q (new_AGEMA_signal_23261) ) ;
    buf_clk new_AGEMA_reg_buffer_10541 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_23265) ) ;
    buf_clk new_AGEMA_reg_buffer_10545 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_23269) ) ;
    buf_clk new_AGEMA_reg_buffer_10549 ( .C (clk), .D (key_s2[121]), .Q (new_AGEMA_signal_23273) ) ;
    buf_clk new_AGEMA_reg_buffer_10553 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_23277) ) ;
    buf_clk new_AGEMA_reg_buffer_10557 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_23281) ) ;
    buf_clk new_AGEMA_reg_buffer_10561 ( .C (clk), .D (key_s2[122]), .Q (new_AGEMA_signal_23285) ) ;
    buf_clk new_AGEMA_reg_buffer_10565 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_23289) ) ;
    buf_clk new_AGEMA_reg_buffer_10569 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_23293) ) ;
    buf_clk new_AGEMA_reg_buffer_10573 ( .C (clk), .D (key_s2[123]), .Q (new_AGEMA_signal_23297) ) ;
    buf_clk new_AGEMA_reg_buffer_10577 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_23301) ) ;
    buf_clk new_AGEMA_reg_buffer_10581 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_23305) ) ;
    buf_clk new_AGEMA_reg_buffer_10585 ( .C (clk), .D (key_s2[124]), .Q (new_AGEMA_signal_23309) ) ;
    buf_clk new_AGEMA_reg_buffer_10589 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_23313) ) ;
    buf_clk new_AGEMA_reg_buffer_10593 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_23317) ) ;
    buf_clk new_AGEMA_reg_buffer_10597 ( .C (clk), .D (key_s2[125]), .Q (new_AGEMA_signal_23321) ) ;
    buf_clk new_AGEMA_reg_buffer_10601 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_23325) ) ;
    buf_clk new_AGEMA_reg_buffer_10605 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_23329) ) ;
    buf_clk new_AGEMA_reg_buffer_10609 ( .C (clk), .D (key_s2[126]), .Q (new_AGEMA_signal_23333) ) ;
    buf_clk new_AGEMA_reg_buffer_10613 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_23337) ) ;
    buf_clk new_AGEMA_reg_buffer_10617 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_23341) ) ;
    buf_clk new_AGEMA_reg_buffer_10621 ( .C (clk), .D (key_s2[127]), .Q (new_AGEMA_signal_23345) ) ;
    buf_clk new_AGEMA_reg_buffer_10625 ( .C (clk), .D (RoundKey[9]), .Q (new_AGEMA_signal_23349) ) ;
    buf_clk new_AGEMA_reg_buffer_10629 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_23353) ) ;
    buf_clk new_AGEMA_reg_buffer_10633 ( .C (clk), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_23357) ) ;
    buf_clk new_AGEMA_reg_buffer_10637 ( .C (clk), .D (RoundKey[8]), .Q (new_AGEMA_signal_23361) ) ;
    buf_clk new_AGEMA_reg_buffer_10641 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_23365) ) ;
    buf_clk new_AGEMA_reg_buffer_10645 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_23369) ) ;
    buf_clk new_AGEMA_reg_buffer_10649 ( .C (clk), .D (RoundKey[7]), .Q (new_AGEMA_signal_23373) ) ;
    buf_clk new_AGEMA_reg_buffer_10653 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_23377) ) ;
    buf_clk new_AGEMA_reg_buffer_10657 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_23381) ) ;
    buf_clk new_AGEMA_reg_buffer_10661 ( .C (clk), .D (RoundKey[6]), .Q (new_AGEMA_signal_23385) ) ;
    buf_clk new_AGEMA_reg_buffer_10665 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_23389) ) ;
    buf_clk new_AGEMA_reg_buffer_10669 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_23393) ) ;
    buf_clk new_AGEMA_reg_buffer_10673 ( .C (clk), .D (RoundKey[5]), .Q (new_AGEMA_signal_23397) ) ;
    buf_clk new_AGEMA_reg_buffer_10677 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_23401) ) ;
    buf_clk new_AGEMA_reg_buffer_10681 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_23405) ) ;
    buf_clk new_AGEMA_reg_buffer_10685 ( .C (clk), .D (RoundKey[4]), .Q (new_AGEMA_signal_23409) ) ;
    buf_clk new_AGEMA_reg_buffer_10689 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_23413) ) ;
    buf_clk new_AGEMA_reg_buffer_10693 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_23417) ) ;
    buf_clk new_AGEMA_reg_buffer_10697 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_23421) ) ;
    buf_clk new_AGEMA_reg_buffer_10701 ( .C (clk), .D (new_AGEMA_signal_4929), .Q (new_AGEMA_signal_23425) ) ;
    buf_clk new_AGEMA_reg_buffer_10705 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_23429) ) ;
    buf_clk new_AGEMA_reg_buffer_10709 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_23433) ) ;
    buf_clk new_AGEMA_reg_buffer_10713 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_23437) ) ;
    buf_clk new_AGEMA_reg_buffer_10717 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_23441) ) ;
    buf_clk new_AGEMA_reg_buffer_10721 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_23445) ) ;
    buf_clk new_AGEMA_reg_buffer_10725 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_23449) ) ;
    buf_clk new_AGEMA_reg_buffer_10729 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_23453) ) ;
    buf_clk new_AGEMA_reg_buffer_10733 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_23457) ) ;
    buf_clk new_AGEMA_reg_buffer_10737 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_23461) ) ;
    buf_clk new_AGEMA_reg_buffer_10741 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_23465) ) ;
    buf_clk new_AGEMA_reg_buffer_10745 ( .C (clk), .D (RoundKey[3]), .Q (new_AGEMA_signal_23469) ) ;
    buf_clk new_AGEMA_reg_buffer_10749 ( .C (clk), .D (new_AGEMA_signal_4917), .Q (new_AGEMA_signal_23473) ) ;
    buf_clk new_AGEMA_reg_buffer_10753 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_23477) ) ;
    buf_clk new_AGEMA_reg_buffer_10757 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_23481) ) ;
    buf_clk new_AGEMA_reg_buffer_10761 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_23485) ) ;
    buf_clk new_AGEMA_reg_buffer_10765 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_23489) ) ;
    buf_clk new_AGEMA_reg_buffer_10769 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_23493) ) ;
    buf_clk new_AGEMA_reg_buffer_10773 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_23497) ) ;
    buf_clk new_AGEMA_reg_buffer_10777 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_23501) ) ;
    buf_clk new_AGEMA_reg_buffer_10781 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_23505) ) ;
    buf_clk new_AGEMA_reg_buffer_10785 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_23509) ) ;
    buf_clk new_AGEMA_reg_buffer_10789 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_23513) ) ;
    buf_clk new_AGEMA_reg_buffer_10793 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_23517) ) ;
    buf_clk new_AGEMA_reg_buffer_10797 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_23521) ) ;
    buf_clk new_AGEMA_reg_buffer_10801 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_23525) ) ;
    buf_clk new_AGEMA_reg_buffer_10805 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_23529) ) ;
    buf_clk new_AGEMA_reg_buffer_10809 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (new_AGEMA_signal_23533) ) ;
    buf_clk new_AGEMA_reg_buffer_10813 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_23537) ) ;
    buf_clk new_AGEMA_reg_buffer_10817 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_23541) ) ;
    buf_clk new_AGEMA_reg_buffer_10821 ( .C (clk), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_23545) ) ;
    buf_clk new_AGEMA_reg_buffer_10825 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_23549) ) ;
    buf_clk new_AGEMA_reg_buffer_10829 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_23553) ) ;
    buf_clk new_AGEMA_reg_buffer_10833 ( .C (clk), .D (new_AGEMA_signal_4893), .Q (new_AGEMA_signal_23557) ) ;
    buf_clk new_AGEMA_reg_buffer_10837 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_23561) ) ;
    buf_clk new_AGEMA_reg_buffer_10841 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_23565) ) ;
    buf_clk new_AGEMA_reg_buffer_10845 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_23569) ) ;
    buf_clk new_AGEMA_reg_buffer_10849 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_23573) ) ;
    buf_clk new_AGEMA_reg_buffer_10853 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_23577) ) ;
    buf_clk new_AGEMA_reg_buffer_10857 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_23581) ) ;
    buf_clk new_AGEMA_reg_buffer_10861 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_23585) ) ;
    buf_clk new_AGEMA_reg_buffer_10865 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_23589) ) ;
    buf_clk new_AGEMA_reg_buffer_10869 ( .C (clk), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_23593) ) ;
    buf_clk new_AGEMA_reg_buffer_10873 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_23597) ) ;
    buf_clk new_AGEMA_reg_buffer_10877 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_23601) ) ;
    buf_clk new_AGEMA_reg_buffer_10881 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_23605) ) ;
    buf_clk new_AGEMA_reg_buffer_10885 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_23609) ) ;
    buf_clk new_AGEMA_reg_buffer_10889 ( .C (clk), .D (RoundKey[31]), .Q (new_AGEMA_signal_23613) ) ;
    buf_clk new_AGEMA_reg_buffer_10893 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_23617) ) ;
    buf_clk new_AGEMA_reg_buffer_10897 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_23621) ) ;
    buf_clk new_AGEMA_reg_buffer_10901 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_23625) ) ;
    buf_clk new_AGEMA_reg_buffer_10905 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_23629) ) ;
    buf_clk new_AGEMA_reg_buffer_10909 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_23633) ) ;
    buf_clk new_AGEMA_reg_buffer_10913 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_23637) ) ;
    buf_clk new_AGEMA_reg_buffer_10917 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_23641) ) ;
    buf_clk new_AGEMA_reg_buffer_10921 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_23645) ) ;
    buf_clk new_AGEMA_reg_buffer_10925 ( .C (clk), .D (RoundKey[30]), .Q (new_AGEMA_signal_23649) ) ;
    buf_clk new_AGEMA_reg_buffer_10929 ( .C (clk), .D (new_AGEMA_signal_4857), .Q (new_AGEMA_signal_23653) ) ;
    buf_clk new_AGEMA_reg_buffer_10933 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_23657) ) ;
    buf_clk new_AGEMA_reg_buffer_10937 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_23661) ) ;
    buf_clk new_AGEMA_reg_buffer_10941 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_23665) ) ;
    buf_clk new_AGEMA_reg_buffer_10945 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_23669) ) ;
    buf_clk new_AGEMA_reg_buffer_10949 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_23673) ) ;
    buf_clk new_AGEMA_reg_buffer_10953 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_23677) ) ;
    buf_clk new_AGEMA_reg_buffer_10957 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_23681) ) ;
    buf_clk new_AGEMA_reg_buffer_10961 ( .C (clk), .D (RoundKey[2]), .Q (new_AGEMA_signal_23685) ) ;
    buf_clk new_AGEMA_reg_buffer_10965 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_23689) ) ;
    buf_clk new_AGEMA_reg_buffer_10969 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_23693) ) ;
    buf_clk new_AGEMA_reg_buffer_10973 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_23697) ) ;
    buf_clk new_AGEMA_reg_buffer_10977 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_23701) ) ;
    buf_clk new_AGEMA_reg_buffer_10981 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_23705) ) ;
    buf_clk new_AGEMA_reg_buffer_10985 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_23709) ) ;
    buf_clk new_AGEMA_reg_buffer_10989 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_23713) ) ;
    buf_clk new_AGEMA_reg_buffer_10993 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_23717) ) ;
    buf_clk new_AGEMA_reg_buffer_10997 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_23721) ) ;
    buf_clk new_AGEMA_reg_buffer_11001 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_23725) ) ;
    buf_clk new_AGEMA_reg_buffer_11005 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_23729) ) ;
    buf_clk new_AGEMA_reg_buffer_11009 ( .C (clk), .D (RoundKey[29]), .Q (new_AGEMA_signal_23733) ) ;
    buf_clk new_AGEMA_reg_buffer_11013 ( .C (clk), .D (new_AGEMA_signal_4845), .Q (new_AGEMA_signal_23737) ) ;
    buf_clk new_AGEMA_reg_buffer_11017 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_23741) ) ;
    buf_clk new_AGEMA_reg_buffer_11021 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_23745) ) ;
    buf_clk new_AGEMA_reg_buffer_11025 ( .C (clk), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_23749) ) ;
    buf_clk new_AGEMA_reg_buffer_11029 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_23753) ) ;
    buf_clk new_AGEMA_reg_buffer_11033 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_23757) ) ;
    buf_clk new_AGEMA_reg_buffer_11037 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_23761) ) ;
    buf_clk new_AGEMA_reg_buffer_11041 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_23765) ) ;
    buf_clk new_AGEMA_reg_buffer_11045 ( .C (clk), .D (RoundKey[28]), .Q (new_AGEMA_signal_23769) ) ;
    buf_clk new_AGEMA_reg_buffer_11049 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_23773) ) ;
    buf_clk new_AGEMA_reg_buffer_11053 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_23777) ) ;
    buf_clk new_AGEMA_reg_buffer_11057 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_23781) ) ;
    buf_clk new_AGEMA_reg_buffer_11061 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_23785) ) ;
    buf_clk new_AGEMA_reg_buffer_11065 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_23789) ) ;
    buf_clk new_AGEMA_reg_buffer_11069 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_23793) ) ;
    buf_clk new_AGEMA_reg_buffer_11073 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_23797) ) ;
    buf_clk new_AGEMA_reg_buffer_11077 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_23801) ) ;
    buf_clk new_AGEMA_reg_buffer_11081 ( .C (clk), .D (RoundKey[27]), .Q (new_AGEMA_signal_23805) ) ;
    buf_clk new_AGEMA_reg_buffer_11085 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_23809) ) ;
    buf_clk new_AGEMA_reg_buffer_11089 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_23813) ) ;
    buf_clk new_AGEMA_reg_buffer_11093 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_23817) ) ;
    buf_clk new_AGEMA_reg_buffer_11097 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_23821) ) ;
    buf_clk new_AGEMA_reg_buffer_11101 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_23825) ) ;
    buf_clk new_AGEMA_reg_buffer_11105 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_23829) ) ;
    buf_clk new_AGEMA_reg_buffer_11109 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_23833) ) ;
    buf_clk new_AGEMA_reg_buffer_11113 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_23837) ) ;
    buf_clk new_AGEMA_reg_buffer_11117 ( .C (clk), .D (RoundKey[26]), .Q (new_AGEMA_signal_23841) ) ;
    buf_clk new_AGEMA_reg_buffer_11121 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_23845) ) ;
    buf_clk new_AGEMA_reg_buffer_11125 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_23849) ) ;
    buf_clk new_AGEMA_reg_buffer_11129 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_23853) ) ;
    buf_clk new_AGEMA_reg_buffer_11133 ( .C (clk), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_23857) ) ;
    buf_clk new_AGEMA_reg_buffer_11137 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_23861) ) ;
    buf_clk new_AGEMA_reg_buffer_11141 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_23865) ) ;
    buf_clk new_AGEMA_reg_buffer_11145 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_23869) ) ;
    buf_clk new_AGEMA_reg_buffer_11149 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_23873) ) ;
    buf_clk new_AGEMA_reg_buffer_11153 ( .C (clk), .D (RoundKey[25]), .Q (new_AGEMA_signal_23877) ) ;
    buf_clk new_AGEMA_reg_buffer_11157 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_23881) ) ;
    buf_clk new_AGEMA_reg_buffer_11161 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_23885) ) ;
    buf_clk new_AGEMA_reg_buffer_11165 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_23889) ) ;
    buf_clk new_AGEMA_reg_buffer_11169 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_23893) ) ;
    buf_clk new_AGEMA_reg_buffer_11173 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_23897) ) ;
    buf_clk new_AGEMA_reg_buffer_11177 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_23901) ) ;
    buf_clk new_AGEMA_reg_buffer_11181 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_23905) ) ;
    buf_clk new_AGEMA_reg_buffer_11185 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_23909) ) ;
    buf_clk new_AGEMA_reg_buffer_11189 ( .C (clk), .D (RoundKey[24]), .Q (new_AGEMA_signal_23913) ) ;
    buf_clk new_AGEMA_reg_buffer_11193 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_23917) ) ;
    buf_clk new_AGEMA_reg_buffer_11197 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_23921) ) ;
    buf_clk new_AGEMA_reg_buffer_11201 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_23925) ) ;
    buf_clk new_AGEMA_reg_buffer_11205 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_23929) ) ;
    buf_clk new_AGEMA_reg_buffer_11209 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_23933) ) ;
    buf_clk new_AGEMA_reg_buffer_11213 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_23937) ) ;
    buf_clk new_AGEMA_reg_buffer_11217 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_23941) ) ;
    buf_clk new_AGEMA_reg_buffer_11221 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_23945) ) ;
    buf_clk new_AGEMA_reg_buffer_11225 ( .C (clk), .D (RoundKey[23]), .Q (new_AGEMA_signal_23949) ) ;
    buf_clk new_AGEMA_reg_buffer_11229 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_23953) ) ;
    buf_clk new_AGEMA_reg_buffer_11233 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_23957) ) ;
    buf_clk new_AGEMA_reg_buffer_11237 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_23961) ) ;
    buf_clk new_AGEMA_reg_buffer_11241 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_23965) ) ;
    buf_clk new_AGEMA_reg_buffer_11245 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_23969) ) ;
    buf_clk new_AGEMA_reg_buffer_11249 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_23973) ) ;
    buf_clk new_AGEMA_reg_buffer_11253 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_23977) ) ;
    buf_clk new_AGEMA_reg_buffer_11257 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_23981) ) ;
    buf_clk new_AGEMA_reg_buffer_11261 ( .C (clk), .D (RoundKey[22]), .Q (new_AGEMA_signal_23985) ) ;
    buf_clk new_AGEMA_reg_buffer_11265 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_23989) ) ;
    buf_clk new_AGEMA_reg_buffer_11269 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_23993) ) ;
    buf_clk new_AGEMA_reg_buffer_11273 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_23997) ) ;
    buf_clk new_AGEMA_reg_buffer_11277 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_24001) ) ;
    buf_clk new_AGEMA_reg_buffer_11281 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_24005) ) ;
    buf_clk new_AGEMA_reg_buffer_11285 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_24009) ) ;
    buf_clk new_AGEMA_reg_buffer_11289 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_24013) ) ;
    buf_clk new_AGEMA_reg_buffer_11293 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_24017) ) ;
    buf_clk new_AGEMA_reg_buffer_11297 ( .C (clk), .D (RoundKey[21]), .Q (new_AGEMA_signal_24021) ) ;
    buf_clk new_AGEMA_reg_buffer_11301 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_24025) ) ;
    buf_clk new_AGEMA_reg_buffer_11305 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_24029) ) ;
    buf_clk new_AGEMA_reg_buffer_11309 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_24033) ) ;
    buf_clk new_AGEMA_reg_buffer_11313 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_24037) ) ;
    buf_clk new_AGEMA_reg_buffer_11317 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_24041) ) ;
    buf_clk new_AGEMA_reg_buffer_11321 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_24045) ) ;
    buf_clk new_AGEMA_reg_buffer_11325 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_24049) ) ;
    buf_clk new_AGEMA_reg_buffer_11329 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_24053) ) ;
    buf_clk new_AGEMA_reg_buffer_11333 ( .C (clk), .D (RoundKey[20]), .Q (new_AGEMA_signal_24057) ) ;
    buf_clk new_AGEMA_reg_buffer_11337 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_24061) ) ;
    buf_clk new_AGEMA_reg_buffer_11341 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_24065) ) ;
    buf_clk new_AGEMA_reg_buffer_11345 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_24069) ) ;
    buf_clk new_AGEMA_reg_buffer_11349 ( .C (clk), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_24073) ) ;
    buf_clk new_AGEMA_reg_buffer_11353 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_24077) ) ;
    buf_clk new_AGEMA_reg_buffer_11357 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_24081) ) ;
    buf_clk new_AGEMA_reg_buffer_11361 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_24085) ) ;
    buf_clk new_AGEMA_reg_buffer_11365 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_24089) ) ;
    buf_clk new_AGEMA_reg_buffer_11369 ( .C (clk), .D (RoundKey[1]), .Q (new_AGEMA_signal_24093) ) ;
    buf_clk new_AGEMA_reg_buffer_11373 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_24097) ) ;
    buf_clk new_AGEMA_reg_buffer_11377 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_24101) ) ;
    buf_clk new_AGEMA_reg_buffer_11381 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_24105) ) ;
    buf_clk new_AGEMA_reg_buffer_11385 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (new_AGEMA_signal_24109) ) ;
    buf_clk new_AGEMA_reg_buffer_11389 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_24113) ) ;
    buf_clk new_AGEMA_reg_buffer_11393 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_24117) ) ;
    buf_clk new_AGEMA_reg_buffer_11397 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_24121) ) ;
    buf_clk new_AGEMA_reg_buffer_11401 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_24125) ) ;
    buf_clk new_AGEMA_reg_buffer_11405 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_24129) ) ;
    buf_clk new_AGEMA_reg_buffer_11409 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_24133) ) ;
    buf_clk new_AGEMA_reg_buffer_11413 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_24137) ) ;
    buf_clk new_AGEMA_reg_buffer_11417 ( .C (clk), .D (RoundKey[19]), .Q (new_AGEMA_signal_24141) ) ;
    buf_clk new_AGEMA_reg_buffer_11421 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_24145) ) ;
    buf_clk new_AGEMA_reg_buffer_11425 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_24149) ) ;
    buf_clk new_AGEMA_reg_buffer_11429 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_24153) ) ;
    buf_clk new_AGEMA_reg_buffer_11433 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_24157) ) ;
    buf_clk new_AGEMA_reg_buffer_11437 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_24161) ) ;
    buf_clk new_AGEMA_reg_buffer_11441 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_24165) ) ;
    buf_clk new_AGEMA_reg_buffer_11445 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_24169) ) ;
    buf_clk new_AGEMA_reg_buffer_11449 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_24173) ) ;
    buf_clk new_AGEMA_reg_buffer_11453 ( .C (clk), .D (RoundKey[18]), .Q (new_AGEMA_signal_24177) ) ;
    buf_clk new_AGEMA_reg_buffer_11457 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_24181) ) ;
    buf_clk new_AGEMA_reg_buffer_11461 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_24185) ) ;
    buf_clk new_AGEMA_reg_buffer_11465 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_24189) ) ;
    buf_clk new_AGEMA_reg_buffer_11469 ( .C (clk), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_24193) ) ;
    buf_clk new_AGEMA_reg_buffer_11473 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_24197) ) ;
    buf_clk new_AGEMA_reg_buffer_11477 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_24201) ) ;
    buf_clk new_AGEMA_reg_buffer_11481 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_24205) ) ;
    buf_clk new_AGEMA_reg_buffer_11485 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_24209) ) ;
    buf_clk new_AGEMA_reg_buffer_11489 ( .C (clk), .D (RoundKey[17]), .Q (new_AGEMA_signal_24213) ) ;
    buf_clk new_AGEMA_reg_buffer_11493 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_24217) ) ;
    buf_clk new_AGEMA_reg_buffer_11497 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_24221) ) ;
    buf_clk new_AGEMA_reg_buffer_11501 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_24225) ) ;
    buf_clk new_AGEMA_reg_buffer_11505 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_24229) ) ;
    buf_clk new_AGEMA_reg_buffer_11509 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_24233) ) ;
    buf_clk new_AGEMA_reg_buffer_11513 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_24237) ) ;
    buf_clk new_AGEMA_reg_buffer_11517 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_24241) ) ;
    buf_clk new_AGEMA_reg_buffer_11521 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_24245) ) ;
    buf_clk new_AGEMA_reg_buffer_11525 ( .C (clk), .D (RoundKey[16]), .Q (new_AGEMA_signal_24249) ) ;
    buf_clk new_AGEMA_reg_buffer_11529 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_24253) ) ;
    buf_clk new_AGEMA_reg_buffer_11533 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_24257) ) ;
    buf_clk new_AGEMA_reg_buffer_11537 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_24261) ) ;
    buf_clk new_AGEMA_reg_buffer_11541 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_24265) ) ;
    buf_clk new_AGEMA_reg_buffer_11545 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_24269) ) ;
    buf_clk new_AGEMA_reg_buffer_11549 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_24273) ) ;
    buf_clk new_AGEMA_reg_buffer_11553 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_24277) ) ;
    buf_clk new_AGEMA_reg_buffer_11557 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_24281) ) ;
    buf_clk new_AGEMA_reg_buffer_11561 ( .C (clk), .D (RoundKey[15]), .Q (new_AGEMA_signal_24285) ) ;
    buf_clk new_AGEMA_reg_buffer_11565 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_24289) ) ;
    buf_clk new_AGEMA_reg_buffer_11569 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_24293) ) ;
    buf_clk new_AGEMA_reg_buffer_11573 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_24297) ) ;
    buf_clk new_AGEMA_reg_buffer_11577 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_24301) ) ;
    buf_clk new_AGEMA_reg_buffer_11581 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_24305) ) ;
    buf_clk new_AGEMA_reg_buffer_11585 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_24309) ) ;
    buf_clk new_AGEMA_reg_buffer_11589 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_24313) ) ;
    buf_clk new_AGEMA_reg_buffer_11593 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_24317) ) ;
    buf_clk new_AGEMA_reg_buffer_11597 ( .C (clk), .D (RoundKey[14]), .Q (new_AGEMA_signal_24321) ) ;
    buf_clk new_AGEMA_reg_buffer_11601 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_24325) ) ;
    buf_clk new_AGEMA_reg_buffer_11605 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_24329) ) ;
    buf_clk new_AGEMA_reg_buffer_11609 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_24333) ) ;
    buf_clk new_AGEMA_reg_buffer_11613 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_24337) ) ;
    buf_clk new_AGEMA_reg_buffer_11617 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_24341) ) ;
    buf_clk new_AGEMA_reg_buffer_11621 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_24345) ) ;
    buf_clk new_AGEMA_reg_buffer_11625 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_24349) ) ;
    buf_clk new_AGEMA_reg_buffer_11629 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_24353) ) ;
    buf_clk new_AGEMA_reg_buffer_11633 ( .C (clk), .D (RoundKey[13]), .Q (new_AGEMA_signal_24357) ) ;
    buf_clk new_AGEMA_reg_buffer_11637 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_24361) ) ;
    buf_clk new_AGEMA_reg_buffer_11641 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_24365) ) ;
    buf_clk new_AGEMA_reg_buffer_11645 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_24369) ) ;
    buf_clk new_AGEMA_reg_buffer_11649 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_24373) ) ;
    buf_clk new_AGEMA_reg_buffer_11653 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_24377) ) ;
    buf_clk new_AGEMA_reg_buffer_11657 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_24381) ) ;
    buf_clk new_AGEMA_reg_buffer_11661 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_24385) ) ;
    buf_clk new_AGEMA_reg_buffer_11665 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_24389) ) ;
    buf_clk new_AGEMA_reg_buffer_11669 ( .C (clk), .D (RoundKey[12]), .Q (new_AGEMA_signal_24393) ) ;
    buf_clk new_AGEMA_reg_buffer_11673 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_24397) ) ;
    buf_clk new_AGEMA_reg_buffer_11677 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_24401) ) ;
    buf_clk new_AGEMA_reg_buffer_11681 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_24405) ) ;
    buf_clk new_AGEMA_reg_buffer_11685 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_24409) ) ;
    buf_clk new_AGEMA_reg_buffer_11689 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_24413) ) ;
    buf_clk new_AGEMA_reg_buffer_11693 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_24417) ) ;
    buf_clk new_AGEMA_reg_buffer_11697 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_24421) ) ;
    buf_clk new_AGEMA_reg_buffer_11701 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_24425) ) ;
    buf_clk new_AGEMA_reg_buffer_11705 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_24429) ) ;
    buf_clk new_AGEMA_reg_buffer_11709 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_24433) ) ;
    buf_clk new_AGEMA_reg_buffer_11713 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_24437) ) ;
    buf_clk new_AGEMA_reg_buffer_11717 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_24441) ) ;
    buf_clk new_AGEMA_reg_buffer_11721 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_24445) ) ;
    buf_clk new_AGEMA_reg_buffer_11725 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_24449) ) ;
    buf_clk new_AGEMA_reg_buffer_11729 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_24453) ) ;
    buf_clk new_AGEMA_reg_buffer_11733 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_24457) ) ;
    buf_clk new_AGEMA_reg_buffer_11737 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_24461) ) ;
    buf_clk new_AGEMA_reg_buffer_11741 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_24465) ) ;
    buf_clk new_AGEMA_reg_buffer_11745 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_24469) ) ;
    buf_clk new_AGEMA_reg_buffer_11749 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_24473) ) ;
    buf_clk new_AGEMA_reg_buffer_11753 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_24477) ) ;
    buf_clk new_AGEMA_reg_buffer_11757 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_24481) ) ;
    buf_clk new_AGEMA_reg_buffer_11761 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_24485) ) ;
    buf_clk new_AGEMA_reg_buffer_11765 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_24489) ) ;
    buf_clk new_AGEMA_reg_buffer_11769 ( .C (clk), .D (new_AGEMA_signal_4701), .Q (new_AGEMA_signal_24493) ) ;
    buf_clk new_AGEMA_reg_buffer_11773 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_24497) ) ;
    buf_clk new_AGEMA_reg_buffer_11777 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_24501) ) ;
    buf_clk new_AGEMA_reg_buffer_11781 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_24505) ) ;
    buf_clk new_AGEMA_reg_buffer_11785 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_24509) ) ;
    buf_clk new_AGEMA_reg_buffer_11789 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_24513) ) ;
    buf_clk new_AGEMA_reg_buffer_11793 ( .C (clk), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_24517) ) ;
    buf_clk new_AGEMA_reg_buffer_11797 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_24521) ) ;
    buf_clk new_AGEMA_reg_buffer_11801 ( .C (clk), .D (RoundKey[11]), .Q (new_AGEMA_signal_24525) ) ;
    buf_clk new_AGEMA_reg_buffer_11805 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_24529) ) ;
    buf_clk new_AGEMA_reg_buffer_11809 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_24533) ) ;
    buf_clk new_AGEMA_reg_buffer_11813 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_24537) ) ;
    buf_clk new_AGEMA_reg_buffer_11817 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_24541) ) ;
    buf_clk new_AGEMA_reg_buffer_11821 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_24545) ) ;
    buf_clk new_AGEMA_reg_buffer_11825 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_24549) ) ;
    buf_clk new_AGEMA_reg_buffer_11829 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_24553) ) ;
    buf_clk new_AGEMA_reg_buffer_11833 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_24557) ) ;
    buf_clk new_AGEMA_reg_buffer_11837 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_24561) ) ;
    buf_clk new_AGEMA_reg_buffer_11841 ( .C (clk), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_24565) ) ;
    buf_clk new_AGEMA_reg_buffer_11845 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_24569) ) ;
    buf_clk new_AGEMA_reg_buffer_11849 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_24573) ) ;
    buf_clk new_AGEMA_reg_buffer_11853 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_24577) ) ;
    buf_clk new_AGEMA_reg_buffer_11857 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_24581) ) ;
    buf_clk new_AGEMA_reg_buffer_11861 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_24585) ) ;
    buf_clk new_AGEMA_reg_buffer_11865 ( .C (clk), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_24589) ) ;
    buf_clk new_AGEMA_reg_buffer_11869 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_24593) ) ;
    buf_clk new_AGEMA_reg_buffer_11873 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_24597) ) ;
    buf_clk new_AGEMA_reg_buffer_11877 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_24601) ) ;
    buf_clk new_AGEMA_reg_buffer_11881 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_24605) ) ;
    buf_clk new_AGEMA_reg_buffer_11885 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_24609) ) ;
    buf_clk new_AGEMA_reg_buffer_11889 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_24613) ) ;
    buf_clk new_AGEMA_reg_buffer_11893 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_24617) ) ;
    buf_clk new_AGEMA_reg_buffer_11897 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_24621) ) ;
    buf_clk new_AGEMA_reg_buffer_11901 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_24625) ) ;
    buf_clk new_AGEMA_reg_buffer_11905 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_24629) ) ;
    buf_clk new_AGEMA_reg_buffer_11909 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_24633) ) ;
    buf_clk new_AGEMA_reg_buffer_11913 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_24637) ) ;
    buf_clk new_AGEMA_reg_buffer_11917 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_24641) ) ;
    buf_clk new_AGEMA_reg_buffer_11921 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_24645) ) ;
    buf_clk new_AGEMA_reg_buffer_11925 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_24649) ) ;
    buf_clk new_AGEMA_reg_buffer_11929 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_24653) ) ;
    buf_clk new_AGEMA_reg_buffer_11933 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_24657) ) ;
    buf_clk new_AGEMA_reg_buffer_11937 ( .C (clk), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_24661) ) ;
    buf_clk new_AGEMA_reg_buffer_11941 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_24665) ) ;
    buf_clk new_AGEMA_reg_buffer_11945 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_24669) ) ;
    buf_clk new_AGEMA_reg_buffer_11949 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_24673) ) ;
    buf_clk new_AGEMA_reg_buffer_11953 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_24677) ) ;
    buf_clk new_AGEMA_reg_buffer_11957 ( .C (clk), .D (RoundKey[10]), .Q (new_AGEMA_signal_24681) ) ;
    buf_clk new_AGEMA_reg_buffer_11961 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_24685) ) ;
    buf_clk new_AGEMA_reg_buffer_11965 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_24689) ) ;
    buf_clk new_AGEMA_reg_buffer_11969 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_24693) ) ;
    buf_clk new_AGEMA_reg_buffer_11973 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_24697) ) ;
    buf_clk new_AGEMA_reg_buffer_11977 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_24701) ) ;
    buf_clk new_AGEMA_reg_buffer_11981 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_24705) ) ;
    buf_clk new_AGEMA_reg_buffer_11985 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_24709) ) ;
    buf_clk new_AGEMA_reg_buffer_11989 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_24713) ) ;
    buf_clk new_AGEMA_reg_buffer_11993 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_24717) ) ;
    buf_clk new_AGEMA_reg_buffer_11997 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_24721) ) ;
    buf_clk new_AGEMA_reg_buffer_12001 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_24725) ) ;
    buf_clk new_AGEMA_reg_buffer_12005 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_24729) ) ;
    buf_clk new_AGEMA_reg_buffer_12009 ( .C (clk), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_24733) ) ;
    buf_clk new_AGEMA_reg_buffer_12013 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_24737) ) ;
    buf_clk new_AGEMA_reg_buffer_12017 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_24741) ) ;
    buf_clk new_AGEMA_reg_buffer_12021 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_24745) ) ;
    buf_clk new_AGEMA_reg_buffer_12025 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_24749) ) ;
    buf_clk new_AGEMA_reg_buffer_12029 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_24753) ) ;
    buf_clk new_AGEMA_reg_buffer_12033 ( .C (clk), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_24757) ) ;
    buf_clk new_AGEMA_reg_buffer_12037 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_24761) ) ;
    buf_clk new_AGEMA_reg_buffer_12041 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_24765) ) ;
    buf_clk new_AGEMA_reg_buffer_12045 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_24769) ) ;
    buf_clk new_AGEMA_reg_buffer_12049 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_24773) ) ;
    buf_clk new_AGEMA_reg_buffer_12053 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_24777) ) ;
    buf_clk new_AGEMA_reg_buffer_12057 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_24781) ) ;
    buf_clk new_AGEMA_reg_buffer_12061 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_24785) ) ;
    buf_clk new_AGEMA_reg_buffer_12065 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_24789) ) ;
    buf_clk new_AGEMA_reg_buffer_12069 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_24793) ) ;
    buf_clk new_AGEMA_reg_buffer_12073 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_24797) ) ;
    buf_clk new_AGEMA_reg_buffer_12077 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_24801) ) ;
    buf_clk new_AGEMA_reg_buffer_12081 ( .C (clk), .D (new_AGEMA_signal_4569), .Q (new_AGEMA_signal_24805) ) ;
    buf_clk new_AGEMA_reg_buffer_12085 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_24809) ) ;
    buf_clk new_AGEMA_reg_buffer_12089 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_24813) ) ;
    buf_clk new_AGEMA_reg_buffer_12093 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_24817) ) ;
    buf_clk new_AGEMA_reg_buffer_12097 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_24821) ) ;
    buf_clk new_AGEMA_reg_buffer_12101 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_24825) ) ;
    buf_clk new_AGEMA_reg_buffer_12105 ( .C (clk), .D (new_AGEMA_signal_4557), .Q (new_AGEMA_signal_24829) ) ;
    buf_clk new_AGEMA_reg_buffer_12109 ( .C (clk), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_24833) ) ;
    buf_clk new_AGEMA_reg_buffer_12113 ( .C (clk), .D (RoundKey[0]), .Q (new_AGEMA_signal_24837) ) ;
    buf_clk new_AGEMA_reg_buffer_12117 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_24841) ) ;
    buf_clk new_AGEMA_reg_buffer_12121 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_24845) ) ;
    buf_clk new_AGEMA_reg_buffer_12125 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_24849) ) ;
    buf_clk new_AGEMA_reg_buffer_12129 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_24853) ) ;
    buf_clk new_AGEMA_reg_buffer_12133 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_24857) ) ;
    buf_clk new_AGEMA_reg_buffer_12137 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_24861) ) ;
    buf_clk new_AGEMA_reg_buffer_12141 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_24865) ) ;
    buf_clk new_AGEMA_reg_buffer_12145 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_24869) ) ;
    buf_clk new_AGEMA_reg_buffer_12149 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_24873) ) ;
    buf_clk new_AGEMA_reg_buffer_12153 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_24877) ) ;
    buf_clk new_AGEMA_reg_buffer_12157 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_24881) ) ;
    buf_clk new_AGEMA_reg_buffer_12161 ( .C (clk), .D (n283), .Q (new_AGEMA_signal_24885) ) ;
    buf_clk new_AGEMA_reg_buffer_12165 ( .C (clk), .D (n285), .Q (new_AGEMA_signal_24889) ) ;
    buf_clk new_AGEMA_reg_buffer_12169 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_24893) ) ;
    buf_clk new_AGEMA_reg_buffer_12173 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_24897) ) ;
    buf_clk new_AGEMA_reg_buffer_12177 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_24901) ) ;
    buf_clk new_AGEMA_reg_buffer_12181 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_24905) ) ;
    buf_clk new_AGEMA_reg_buffer_12185 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_24909) ) ;
    buf_clk new_AGEMA_reg_buffer_12189 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_24913) ) ;
    buf_clk new_AGEMA_reg_buffer_12193 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_24917) ) ;
    buf_clk new_AGEMA_reg_buffer_12196 ( .C (clk), .D (new_AGEMA_signal_5717), .Q (new_AGEMA_signal_24920) ) ;
    buf_clk new_AGEMA_reg_buffer_12199 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_24923) ) ;
    buf_clk new_AGEMA_reg_buffer_12202 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_24926) ) ;
    buf_clk new_AGEMA_reg_buffer_12205 ( .C (clk), .D (new_AGEMA_signal_6037), .Q (new_AGEMA_signal_24929) ) ;
    buf_clk new_AGEMA_reg_buffer_12208 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_24932) ) ;
    buf_clk new_AGEMA_reg_buffer_12211 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_24935) ) ;
    buf_clk new_AGEMA_reg_buffer_12214 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_24938) ) ;
    buf_clk new_AGEMA_reg_buffer_12217 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_24941) ) ;
    buf_clk new_AGEMA_reg_buffer_12220 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_24944) ) ;
    buf_clk new_AGEMA_reg_buffer_12223 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_24947) ) ;
    buf_clk new_AGEMA_reg_buffer_12226 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_24950) ) ;
    buf_clk new_AGEMA_reg_buffer_12229 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_24953) ) ;
    buf_clk new_AGEMA_reg_buffer_12232 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_24956) ) ;
    buf_clk new_AGEMA_reg_buffer_12235 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_24959) ) ;
    buf_clk new_AGEMA_reg_buffer_12238 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_24962) ) ;
    buf_clk new_AGEMA_reg_buffer_12241 ( .C (clk), .D (new_AGEMA_signal_5723), .Q (new_AGEMA_signal_24965) ) ;
    buf_clk new_AGEMA_reg_buffer_12244 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_24968) ) ;
    buf_clk new_AGEMA_reg_buffer_12247 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_24971) ) ;
    buf_clk new_AGEMA_reg_buffer_12250 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_24974) ) ;
    buf_clk new_AGEMA_reg_buffer_12253 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_24977) ) ;
    buf_clk new_AGEMA_reg_buffer_12256 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_24980) ) ;
    buf_clk new_AGEMA_reg_buffer_12259 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_24983) ) ;
    buf_clk new_AGEMA_reg_buffer_12262 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_24986) ) ;
    buf_clk new_AGEMA_reg_buffer_12265 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_24989) ) ;
    buf_clk new_AGEMA_reg_buffer_12268 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_24992) ) ;
    buf_clk new_AGEMA_reg_buffer_12271 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_24995) ) ;
    buf_clk new_AGEMA_reg_buffer_12274 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_24998) ) ;
    buf_clk new_AGEMA_reg_buffer_12277 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_25001) ) ;
    buf_clk new_AGEMA_reg_buffer_12280 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_25004) ) ;
    buf_clk new_AGEMA_reg_buffer_12283 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_25007) ) ;
    buf_clk new_AGEMA_reg_buffer_12286 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_25010) ) ;
    buf_clk new_AGEMA_reg_buffer_12289 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_25013) ) ;
    buf_clk new_AGEMA_reg_buffer_12292 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_25016) ) ;
    buf_clk new_AGEMA_reg_buffer_12295 ( .C (clk), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_25019) ) ;
    buf_clk new_AGEMA_reg_buffer_12298 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_25022) ) ;
    buf_clk new_AGEMA_reg_buffer_12301 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_25025) ) ;
    buf_clk new_AGEMA_reg_buffer_12304 ( .C (clk), .D (new_AGEMA_signal_5729), .Q (new_AGEMA_signal_25028) ) ;
    buf_clk new_AGEMA_reg_buffer_12307 ( .C (clk), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_25031) ) ;
    buf_clk new_AGEMA_reg_buffer_12310 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_25034) ) ;
    buf_clk new_AGEMA_reg_buffer_12313 ( .C (clk), .D (new_AGEMA_signal_6045), .Q (new_AGEMA_signal_25037) ) ;
    buf_clk new_AGEMA_reg_buffer_12316 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_25040) ) ;
    buf_clk new_AGEMA_reg_buffer_12319 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_25043) ) ;
    buf_clk new_AGEMA_reg_buffer_12322 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_25046) ) ;
    buf_clk new_AGEMA_reg_buffer_12325 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_25049) ) ;
    buf_clk new_AGEMA_reg_buffer_12328 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_25052) ) ;
    buf_clk new_AGEMA_reg_buffer_12331 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_25055) ) ;
    buf_clk new_AGEMA_reg_buffer_12334 ( .C (clk), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_25058) ) ;
    buf_clk new_AGEMA_reg_buffer_12337 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_25061) ) ;
    buf_clk new_AGEMA_reg_buffer_12340 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_25064) ) ;
    buf_clk new_AGEMA_reg_buffer_12343 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_25067) ) ;
    buf_clk new_AGEMA_reg_buffer_12346 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_25070) ) ;
    buf_clk new_AGEMA_reg_buffer_12349 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_25073) ) ;
    buf_clk new_AGEMA_reg_buffer_12352 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_25076) ) ;
    buf_clk new_AGEMA_reg_buffer_12355 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_25079) ) ;
    buf_clk new_AGEMA_reg_buffer_12358 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_25082) ) ;
    buf_clk new_AGEMA_reg_buffer_12361 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_25085) ) ;
    buf_clk new_AGEMA_reg_buffer_12364 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_25088) ) ;
    buf_clk new_AGEMA_reg_buffer_12367 ( .C (clk), .D (new_AGEMA_signal_5741), .Q (new_AGEMA_signal_25091) ) ;
    buf_clk new_AGEMA_reg_buffer_12370 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_25094) ) ;
    buf_clk new_AGEMA_reg_buffer_12373 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_25097) ) ;
    buf_clk new_AGEMA_reg_buffer_12376 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_25100) ) ;
    buf_clk new_AGEMA_reg_buffer_12379 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_25103) ) ;
    buf_clk new_AGEMA_reg_buffer_12382 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_25106) ) ;
    buf_clk new_AGEMA_reg_buffer_12385 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_25109) ) ;
    buf_clk new_AGEMA_reg_buffer_12388 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_25112) ) ;
    buf_clk new_AGEMA_reg_buffer_12391 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_25115) ) ;
    buf_clk new_AGEMA_reg_buffer_12394 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_25118) ) ;
    buf_clk new_AGEMA_reg_buffer_12397 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_25121) ) ;
    buf_clk new_AGEMA_reg_buffer_12400 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_25124) ) ;
    buf_clk new_AGEMA_reg_buffer_12403 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_25127) ) ;
    buf_clk new_AGEMA_reg_buffer_12406 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_25130) ) ;
    buf_clk new_AGEMA_reg_buffer_12409 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_25133) ) ;
    buf_clk new_AGEMA_reg_buffer_12412 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_25136) ) ;
    buf_clk new_AGEMA_reg_buffer_12415 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_25139) ) ;
    buf_clk new_AGEMA_reg_buffer_12418 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_25142) ) ;
    buf_clk new_AGEMA_reg_buffer_12421 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_25145) ) ;
    buf_clk new_AGEMA_reg_buffer_12424 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_25148) ) ;
    buf_clk new_AGEMA_reg_buffer_12427 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_25151) ) ;
    buf_clk new_AGEMA_reg_buffer_12430 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_25154) ) ;
    buf_clk new_AGEMA_reg_buffer_12433 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_25157) ) ;
    buf_clk new_AGEMA_reg_buffer_12436 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_25160) ) ;
    buf_clk new_AGEMA_reg_buffer_12439 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_25163) ) ;
    buf_clk new_AGEMA_reg_buffer_12442 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_25166) ) ;
    buf_clk new_AGEMA_reg_buffer_12445 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_25169) ) ;
    buf_clk new_AGEMA_reg_buffer_12448 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_25172) ) ;
    buf_clk new_AGEMA_reg_buffer_12451 ( .C (clk), .D (new_AGEMA_signal_5342), .Q (new_AGEMA_signal_25175) ) ;
    buf_clk new_AGEMA_reg_buffer_12454 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_25178) ) ;
    buf_clk new_AGEMA_reg_buffer_12457 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_25181) ) ;
    buf_clk new_AGEMA_reg_buffer_12460 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_25184) ) ;
    buf_clk new_AGEMA_reg_buffer_12463 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_25187) ) ;
    buf_clk new_AGEMA_reg_buffer_12466 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_25190) ) ;
    buf_clk new_AGEMA_reg_buffer_12469 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_25193) ) ;
    buf_clk new_AGEMA_reg_buffer_12472 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_25196) ) ;
    buf_clk new_AGEMA_reg_buffer_12475 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_25199) ) ;
    buf_clk new_AGEMA_reg_buffer_12478 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_25202) ) ;
    buf_clk new_AGEMA_reg_buffer_12481 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_25205) ) ;
    buf_clk new_AGEMA_reg_buffer_12484 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_25208) ) ;
    buf_clk new_AGEMA_reg_buffer_12487 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_25211) ) ;
    buf_clk new_AGEMA_reg_buffer_12490 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_25214) ) ;
    buf_clk new_AGEMA_reg_buffer_12493 ( .C (clk), .D (new_AGEMA_signal_5339), .Q (new_AGEMA_signal_25217) ) ;
    buf_clk new_AGEMA_reg_buffer_12496 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_25220) ) ;
    buf_clk new_AGEMA_reg_buffer_12499 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_25223) ) ;
    buf_clk new_AGEMA_reg_buffer_12502 ( .C (clk), .D (new_AGEMA_signal_5749), .Q (new_AGEMA_signal_25226) ) ;
    buf_clk new_AGEMA_reg_buffer_12505 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_25229) ) ;
    buf_clk new_AGEMA_reg_buffer_12508 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_25232) ) ;
    buf_clk new_AGEMA_reg_buffer_12511 ( .C (clk), .D (new_AGEMA_signal_6089), .Q (new_AGEMA_signal_25235) ) ;
    buf_clk new_AGEMA_reg_buffer_12514 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_25238) ) ;
    buf_clk new_AGEMA_reg_buffer_12517 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_25241) ) ;
    buf_clk new_AGEMA_reg_buffer_12520 ( .C (clk), .D (new_AGEMA_signal_5757), .Q (new_AGEMA_signal_25244) ) ;
    buf_clk new_AGEMA_reg_buffer_12523 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_25247) ) ;
    buf_clk new_AGEMA_reg_buffer_12526 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_25250) ) ;
    buf_clk new_AGEMA_reg_buffer_12529 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_25253) ) ;
    buf_clk new_AGEMA_reg_buffer_12532 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_25256) ) ;
    buf_clk new_AGEMA_reg_buffer_12535 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_25259) ) ;
    buf_clk new_AGEMA_reg_buffer_12538 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_25262) ) ;
    buf_clk new_AGEMA_reg_buffer_12541 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_25265) ) ;
    buf_clk new_AGEMA_reg_buffer_12544 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_25268) ) ;
    buf_clk new_AGEMA_reg_buffer_12547 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_25271) ) ;
    buf_clk new_AGEMA_reg_buffer_12550 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_25274) ) ;
    buf_clk new_AGEMA_reg_buffer_12553 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_25277) ) ;
    buf_clk new_AGEMA_reg_buffer_12556 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_25280) ) ;
    buf_clk new_AGEMA_reg_buffer_12559 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_25283) ) ;
    buf_clk new_AGEMA_reg_buffer_12562 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_25286) ) ;
    buf_clk new_AGEMA_reg_buffer_12565 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_25289) ) ;
    buf_clk new_AGEMA_reg_buffer_12568 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_25292) ) ;
    buf_clk new_AGEMA_reg_buffer_12571 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_25295) ) ;
    buf_clk new_AGEMA_reg_buffer_12574 ( .C (clk), .D (new_AGEMA_signal_5753), .Q (new_AGEMA_signal_25298) ) ;
    buf_clk new_AGEMA_reg_buffer_12577 ( .C (clk), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_25301) ) ;
    buf_clk new_AGEMA_reg_buffer_12580 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_25304) ) ;
    buf_clk new_AGEMA_reg_buffer_12583 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_25307) ) ;
    buf_clk new_AGEMA_reg_buffer_12586 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_25310) ) ;
    buf_clk new_AGEMA_reg_buffer_12589 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_25313) ) ;
    buf_clk new_AGEMA_reg_buffer_12592 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_25316) ) ;
    buf_clk new_AGEMA_reg_buffer_12595 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_25319) ) ;
    buf_clk new_AGEMA_reg_buffer_12598 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_25322) ) ;
    buf_clk new_AGEMA_reg_buffer_12601 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_25325) ) ;
    buf_clk new_AGEMA_reg_buffer_12604 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_25328) ) ;
    buf_clk new_AGEMA_reg_buffer_12607 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_25331) ) ;
    buf_clk new_AGEMA_reg_buffer_12610 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_25334) ) ;
    buf_clk new_AGEMA_reg_buffer_12613 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_25337) ) ;
    buf_clk new_AGEMA_reg_buffer_12616 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_25340) ) ;
    buf_clk new_AGEMA_reg_buffer_12619 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_25343) ) ;
    buf_clk new_AGEMA_reg_buffer_12622 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_25346) ) ;
    buf_clk new_AGEMA_reg_buffer_12625 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_25349) ) ;
    buf_clk new_AGEMA_reg_buffer_12628 ( .C (clk), .D (new_AGEMA_signal_5357), .Q (new_AGEMA_signal_25352) ) ;
    buf_clk new_AGEMA_reg_buffer_12631 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_25355) ) ;
    buf_clk new_AGEMA_reg_buffer_12634 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_25358) ) ;
    buf_clk new_AGEMA_reg_buffer_12637 ( .C (clk), .D (new_AGEMA_signal_5363), .Q (new_AGEMA_signal_25361) ) ;
    buf_clk new_AGEMA_reg_buffer_12640 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_25364) ) ;
    buf_clk new_AGEMA_reg_buffer_12643 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_25367) ) ;
    buf_clk new_AGEMA_reg_buffer_12646 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_25370) ) ;
    buf_clk new_AGEMA_reg_buffer_12649 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_25373) ) ;
    buf_clk new_AGEMA_reg_buffer_12652 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_25376) ) ;
    buf_clk new_AGEMA_reg_buffer_12655 ( .C (clk), .D (new_AGEMA_signal_5765), .Q (new_AGEMA_signal_25379) ) ;
    buf_clk new_AGEMA_reg_buffer_12658 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_25382) ) ;
    buf_clk new_AGEMA_reg_buffer_12661 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_25385) ) ;
    buf_clk new_AGEMA_reg_buffer_12664 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_25388) ) ;
    buf_clk new_AGEMA_reg_buffer_12667 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_25391) ) ;
    buf_clk new_AGEMA_reg_buffer_12670 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_25394) ) ;
    buf_clk new_AGEMA_reg_buffer_12673 ( .C (clk), .D (new_AGEMA_signal_5773), .Q (new_AGEMA_signal_25397) ) ;
    buf_clk new_AGEMA_reg_buffer_12676 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_25400) ) ;
    buf_clk new_AGEMA_reg_buffer_12679 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_25403) ) ;
    buf_clk new_AGEMA_reg_buffer_12682 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_25406) ) ;
    buf_clk new_AGEMA_reg_buffer_12685 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_25409) ) ;
    buf_clk new_AGEMA_reg_buffer_12688 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_25412) ) ;
    buf_clk new_AGEMA_reg_buffer_12691 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_25415) ) ;
    buf_clk new_AGEMA_reg_buffer_12694 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_25418) ) ;
    buf_clk new_AGEMA_reg_buffer_12697 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_25421) ) ;
    buf_clk new_AGEMA_reg_buffer_12700 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_25424) ) ;
    buf_clk new_AGEMA_reg_buffer_12703 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_25427) ) ;
    buf_clk new_AGEMA_reg_buffer_12706 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_25430) ) ;
    buf_clk new_AGEMA_reg_buffer_12709 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_25433) ) ;
    buf_clk new_AGEMA_reg_buffer_12712 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_25436) ) ;
    buf_clk new_AGEMA_reg_buffer_12715 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_25439) ) ;
    buf_clk new_AGEMA_reg_buffer_12718 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_25442) ) ;
    buf_clk new_AGEMA_reg_buffer_12721 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_25445) ) ;
    buf_clk new_AGEMA_reg_buffer_12724 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_25448) ) ;
    buf_clk new_AGEMA_reg_buffer_12727 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_25451) ) ;
    buf_clk new_AGEMA_reg_buffer_12730 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_25454) ) ;
    buf_clk new_AGEMA_reg_buffer_12733 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_25457) ) ;
    buf_clk new_AGEMA_reg_buffer_12736 ( .C (clk), .D (new_AGEMA_signal_6125), .Q (new_AGEMA_signal_25460) ) ;
    buf_clk new_AGEMA_reg_buffer_12739 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_25463) ) ;
    buf_clk new_AGEMA_reg_buffer_12742 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_25466) ) ;
    buf_clk new_AGEMA_reg_buffer_12745 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_25469) ) ;
    buf_clk new_AGEMA_reg_buffer_12748 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_25472) ) ;
    buf_clk new_AGEMA_reg_buffer_12751 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_25475) ) ;
    buf_clk new_AGEMA_reg_buffer_12754 ( .C (clk), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_25478) ) ;
    buf_clk new_AGEMA_reg_buffer_12757 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_25481) ) ;
    buf_clk new_AGEMA_reg_buffer_12760 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_25484) ) ;
    buf_clk new_AGEMA_reg_buffer_12763 ( .C (clk), .D (new_AGEMA_signal_5777), .Q (new_AGEMA_signal_25487) ) ;
    buf_clk new_AGEMA_reg_buffer_12766 ( .C (clk), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_25490) ) ;
    buf_clk new_AGEMA_reg_buffer_12769 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_25493) ) ;
    buf_clk new_AGEMA_reg_buffer_12772 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_25496) ) ;
    buf_clk new_AGEMA_reg_buffer_12775 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_25499) ) ;
    buf_clk new_AGEMA_reg_buffer_12778 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_25502) ) ;
    buf_clk new_AGEMA_reg_buffer_12781 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_25505) ) ;
    buf_clk new_AGEMA_reg_buffer_12784 ( .C (clk), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_25508) ) ;
    buf_clk new_AGEMA_reg_buffer_12787 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_25511) ) ;
    buf_clk new_AGEMA_reg_buffer_12790 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_25514) ) ;
    buf_clk new_AGEMA_reg_buffer_12793 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_25517) ) ;
    buf_clk new_AGEMA_reg_buffer_12796 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_25520) ) ;
    buf_clk new_AGEMA_reg_buffer_12799 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_25523) ) ;
    buf_clk new_AGEMA_reg_buffer_12802 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_25526) ) ;
    buf_clk new_AGEMA_reg_buffer_12805 ( .C (clk), .D (RoundCounterIns_N7), .Q (new_AGEMA_signal_25529) ) ;
    buf_clk new_AGEMA_reg_buffer_12809 ( .C (clk), .D (RoundCounterIns_N8), .Q (new_AGEMA_signal_25533) ) ;
    buf_clk new_AGEMA_reg_buffer_12813 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_25537) ) ;
    buf_clk new_AGEMA_reg_buffer_12817 ( .C (clk), .D (RoundCounterIns_N10), .Q (new_AGEMA_signal_25541) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_17175, new_AGEMA_signal_17174, new_AGEMA_signal_17173}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_17178, new_AGEMA_signal_17177, new_AGEMA_signal_17176}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_17181, new_AGEMA_signal_17180, new_AGEMA_signal_17179}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_17184, new_AGEMA_signal_17183, new_AGEMA_signal_17182}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_17187, new_AGEMA_signal_17186, new_AGEMA_signal_17185}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_17190, new_AGEMA_signal_17189, new_AGEMA_signal_17188}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_17193, new_AGEMA_signal_17192, new_AGEMA_signal_17191}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_17196, new_AGEMA_signal_17195, new_AGEMA_signal_17194}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7696, new_AGEMA_signal_7695, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_17199, new_AGEMA_signal_17198, new_AGEMA_signal_17197}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_17202, new_AGEMA_signal_17201, new_AGEMA_signal_17200}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_17205, new_AGEMA_signal_17204, new_AGEMA_signal_17203}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_17208, new_AGEMA_signal_17207, new_AGEMA_signal_17206}), .b ({new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_17211, new_AGEMA_signal_17210, new_AGEMA_signal_17209}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_17214, new_AGEMA_signal_17213, new_AGEMA_signal_17212}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_17217, new_AGEMA_signal_17216, new_AGEMA_signal_17215}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7516, new_AGEMA_signal_7515, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_17220, new_AGEMA_signal_17219, new_AGEMA_signal_17218}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_17223, new_AGEMA_signal_17222, new_AGEMA_signal_17221}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_17226, new_AGEMA_signal_17225, new_AGEMA_signal_17224}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_17229, new_AGEMA_signal_17228, new_AGEMA_signal_17227}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_17232, new_AGEMA_signal_17231, new_AGEMA_signal_17230}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_7726, new_AGEMA_signal_7725, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_17235, new_AGEMA_signal_17234, new_AGEMA_signal_17233}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_17238, new_AGEMA_signal_17237, new_AGEMA_signal_17236}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_17241, new_AGEMA_signal_17240, new_AGEMA_signal_17239}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_17244, new_AGEMA_signal_17243, new_AGEMA_signal_17242}), .b ({new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_17247, new_AGEMA_signal_17246, new_AGEMA_signal_17245}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_17250, new_AGEMA_signal_17249, new_AGEMA_signal_17248}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_17253, new_AGEMA_signal_17252, new_AGEMA_signal_17251}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7546, new_AGEMA_signal_7545, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_17256, new_AGEMA_signal_17255, new_AGEMA_signal_17254}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_17259, new_AGEMA_signal_17258, new_AGEMA_signal_17257}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_17262, new_AGEMA_signal_17261, new_AGEMA_signal_17260}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_17265, new_AGEMA_signal_17264, new_AGEMA_signal_17263}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_17268, new_AGEMA_signal_17267, new_AGEMA_signal_17266}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_7756, new_AGEMA_signal_7755, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_17271, new_AGEMA_signal_17270, new_AGEMA_signal_17269}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_17274, new_AGEMA_signal_17273, new_AGEMA_signal_17272}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7562, new_AGEMA_signal_7561, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_17277, new_AGEMA_signal_17276, new_AGEMA_signal_17275}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_17280, new_AGEMA_signal_17279, new_AGEMA_signal_17278}), .b ({new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_17283, new_AGEMA_signal_17282, new_AGEMA_signal_17281}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_17286, new_AGEMA_signal_17285, new_AGEMA_signal_17284}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_7574, new_AGEMA_signal_7573, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_17289, new_AGEMA_signal_17288, new_AGEMA_signal_17287}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7576, new_AGEMA_signal_7575, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_17292, new_AGEMA_signal_17291, new_AGEMA_signal_17290}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_17295, new_AGEMA_signal_17294, new_AGEMA_signal_17293}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7580, new_AGEMA_signal_7579, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_17298, new_AGEMA_signal_17297, new_AGEMA_signal_17296}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_17301, new_AGEMA_signal_17300, new_AGEMA_signal_17299}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7586, new_AGEMA_signal_7585, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_17304, new_AGEMA_signal_17303, new_AGEMA_signal_17302}), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_7786, new_AGEMA_signal_7785, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_17307, new_AGEMA_signal_17306, new_AGEMA_signal_17305}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_17310, new_AGEMA_signal_17309, new_AGEMA_signal_17308}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7592, new_AGEMA_signal_7591, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_17313, new_AGEMA_signal_17312, new_AGEMA_signal_17311}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_17316, new_AGEMA_signal_17315, new_AGEMA_signal_17314}), .b ({new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_17319, new_AGEMA_signal_17318, new_AGEMA_signal_17317}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_17322, new_AGEMA_signal_17321, new_AGEMA_signal_17320}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_7604, new_AGEMA_signal_7603, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_17325, new_AGEMA_signal_17324, new_AGEMA_signal_17323}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7606, new_AGEMA_signal_7605, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_17328, new_AGEMA_signal_17327, new_AGEMA_signal_17326}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_17331, new_AGEMA_signal_17330, new_AGEMA_signal_17329}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7610, new_AGEMA_signal_7609, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_17334, new_AGEMA_signal_17333, new_AGEMA_signal_17332}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_17337, new_AGEMA_signal_17336, new_AGEMA_signal_17335}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7616, new_AGEMA_signal_7615, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_17340, new_AGEMA_signal_17339, new_AGEMA_signal_17338}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_7816, new_AGEMA_signal_7815, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_17343, new_AGEMA_signal_17342, new_AGEMA_signal_17341}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_17346, new_AGEMA_signal_17345, new_AGEMA_signal_17344}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7622, new_AGEMA_signal_7621, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_17349, new_AGEMA_signal_17348, new_AGEMA_signal_17347}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_17352, new_AGEMA_signal_17351, new_AGEMA_signal_17350}), .b ({new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_17355, new_AGEMA_signal_17354, new_AGEMA_signal_17353}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_17358, new_AGEMA_signal_17357, new_AGEMA_signal_17356}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_7634, new_AGEMA_signal_7633, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_17361, new_AGEMA_signal_17360, new_AGEMA_signal_17359}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7636, new_AGEMA_signal_7635, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_17364, new_AGEMA_signal_17363, new_AGEMA_signal_17362}), .b ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_17367, new_AGEMA_signal_17366, new_AGEMA_signal_17365}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_17370, new_AGEMA_signal_17369, new_AGEMA_signal_17368}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7442, new_AGEMA_signal_7441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_17373, new_AGEMA_signal_17372, new_AGEMA_signal_17371}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_17376, new_AGEMA_signal_17375, new_AGEMA_signal_17374}), .b ({new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_17379, new_AGEMA_signal_17378, new_AGEMA_signal_17377}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_17382, new_AGEMA_signal_17381, new_AGEMA_signal_17380}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_7454, new_AGEMA_signal_7453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_17385, new_AGEMA_signal_17384, new_AGEMA_signal_17383}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7456, new_AGEMA_signal_7455, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_17388, new_AGEMA_signal_17387, new_AGEMA_signal_17386}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_17391, new_AGEMA_signal_17390, new_AGEMA_signal_17389}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7460, new_AGEMA_signal_7459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_17394, new_AGEMA_signal_17393, new_AGEMA_signal_17392}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_17397, new_AGEMA_signal_17396, new_AGEMA_signal_17395}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7466, new_AGEMA_signal_7465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_17400, new_AGEMA_signal_17399, new_AGEMA_signal_17398}), .b ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_7666, new_AGEMA_signal_7665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_17403, new_AGEMA_signal_17402, new_AGEMA_signal_17401}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_17406, new_AGEMA_signal_17405, new_AGEMA_signal_17404}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7472, new_AGEMA_signal_7471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_17409, new_AGEMA_signal_17408, new_AGEMA_signal_17407}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_17412, new_AGEMA_signal_17411, new_AGEMA_signal_17410}), .b ({new_AGEMA_signal_7304, new_AGEMA_signal_7303, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_7676, new_AGEMA_signal_7675, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_17173) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_7153), .Q (new_AGEMA_signal_17174) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_7154), .Q (new_AGEMA_signal_17175) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_17176) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_7309), .Q (new_AGEMA_signal_17177) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_7310), .Q (new_AGEMA_signal_17178) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_17179) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_7313), .Q (new_AGEMA_signal_17180) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (new_AGEMA_signal_7314), .Q (new_AGEMA_signal_17181) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_17182) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_7477), .Q (new_AGEMA_signal_17183) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_17184) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_17185) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_7161), .Q (new_AGEMA_signal_17186) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_7162), .Q (new_AGEMA_signal_17187) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_17188) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (new_AGEMA_signal_7317), .Q (new_AGEMA_signal_17189) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_7318), .Q (new_AGEMA_signal_17190) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_17191) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_7321), .Q (new_AGEMA_signal_17192) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_7322), .Q (new_AGEMA_signal_17193) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_17194) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_17195) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_17196) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_17197) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_7169), .Q (new_AGEMA_signal_17198) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_7170), .Q (new_AGEMA_signal_17199) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_17200) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (new_AGEMA_signal_7325), .Q (new_AGEMA_signal_17201) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_7326), .Q (new_AGEMA_signal_17202) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_17203) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_7329), .Q (new_AGEMA_signal_17204) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_17205) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_17206) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_7497), .Q (new_AGEMA_signal_17207) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_17208) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_17209) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_7177), .Q (new_AGEMA_signal_17210) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_7178), .Q (new_AGEMA_signal_17211) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_17212) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (new_AGEMA_signal_7333), .Q (new_AGEMA_signal_17213) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_17214) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_17215) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_7337), .Q (new_AGEMA_signal_17216) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_17217) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_17218) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_17219) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_17220) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M21), .Q (new_AGEMA_signal_17221) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_17222) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_17223) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M23), .Q (new_AGEMA_signal_17224) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_7341), .Q (new_AGEMA_signal_17225) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_17226) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M27), .Q (new_AGEMA_signal_17227) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_7345), .Q (new_AGEMA_signal_17228) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_17229) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M24), .Q (new_AGEMA_signal_17230) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_7517), .Q (new_AGEMA_signal_17231) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_17232) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M21), .Q (new_AGEMA_signal_17233) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7193), .Q (new_AGEMA_signal_17234) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_7194), .Q (new_AGEMA_signal_17235) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M23), .Q (new_AGEMA_signal_17236) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (new_AGEMA_signal_7349), .Q (new_AGEMA_signal_17237) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_7350), .Q (new_AGEMA_signal_17238) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M27), .Q (new_AGEMA_signal_17239) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_7353), .Q (new_AGEMA_signal_17240) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (new_AGEMA_signal_7354), .Q (new_AGEMA_signal_17241) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M24), .Q (new_AGEMA_signal_17242) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_17243) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_17244) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M21), .Q (new_AGEMA_signal_17245) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7201), .Q (new_AGEMA_signal_17246) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_7202), .Q (new_AGEMA_signal_17247) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M23), .Q (new_AGEMA_signal_17248) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (new_AGEMA_signal_7357), .Q (new_AGEMA_signal_17249) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7358), .Q (new_AGEMA_signal_17250) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M27), .Q (new_AGEMA_signal_17251) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_7361), .Q (new_AGEMA_signal_17252) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (new_AGEMA_signal_7362), .Q (new_AGEMA_signal_17253) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M24), .Q (new_AGEMA_signal_17254) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_7537), .Q (new_AGEMA_signal_17255) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_17256) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M21), .Q (new_AGEMA_signal_17257) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_7209), .Q (new_AGEMA_signal_17258) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_7210), .Q (new_AGEMA_signal_17259) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M23), .Q (new_AGEMA_signal_17260) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_7365), .Q (new_AGEMA_signal_17261) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_17262) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M27), .Q (new_AGEMA_signal_17263) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_7369), .Q (new_AGEMA_signal_17264) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_17265) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M24), .Q (new_AGEMA_signal_17266) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_7547), .Q (new_AGEMA_signal_17267) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_17268) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M21), .Q (new_AGEMA_signal_17269) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_7217), .Q (new_AGEMA_signal_17270) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_7218), .Q (new_AGEMA_signal_17271) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M23), .Q (new_AGEMA_signal_17272) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_7373), .Q (new_AGEMA_signal_17273) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_17274) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M27), .Q (new_AGEMA_signal_17275) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_7377), .Q (new_AGEMA_signal_17276) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_17277) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M24), .Q (new_AGEMA_signal_17278) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_7557), .Q (new_AGEMA_signal_17279) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_7558), .Q (new_AGEMA_signal_17280) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M21), .Q (new_AGEMA_signal_17281) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_7225), .Q (new_AGEMA_signal_17282) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_17283) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M23), .Q (new_AGEMA_signal_17284) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_7381), .Q (new_AGEMA_signal_17285) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_17286) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M27), .Q (new_AGEMA_signal_17287) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_7385), .Q (new_AGEMA_signal_17288) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_17289) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M24), .Q (new_AGEMA_signal_17290) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_17291) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_17292) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M21), .Q (new_AGEMA_signal_17293) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_7233), .Q (new_AGEMA_signal_17294) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_7234), .Q (new_AGEMA_signal_17295) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M23), .Q (new_AGEMA_signal_17296) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_7389), .Q (new_AGEMA_signal_17297) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_7390), .Q (new_AGEMA_signal_17298) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M27), .Q (new_AGEMA_signal_17299) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_7393), .Q (new_AGEMA_signal_17300) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (new_AGEMA_signal_7394), .Q (new_AGEMA_signal_17301) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M24), .Q (new_AGEMA_signal_17302) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_7577), .Q (new_AGEMA_signal_17303) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_7578), .Q (new_AGEMA_signal_17304) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M21), .Q (new_AGEMA_signal_17305) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_7241), .Q (new_AGEMA_signal_17306) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_7242), .Q (new_AGEMA_signal_17307) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M23), .Q (new_AGEMA_signal_17308) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_7397), .Q (new_AGEMA_signal_17309) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_7398), .Q (new_AGEMA_signal_17310) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M27), .Q (new_AGEMA_signal_17311) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_7401), .Q (new_AGEMA_signal_17312) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_7402), .Q (new_AGEMA_signal_17313) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M24), .Q (new_AGEMA_signal_17314) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_7587), .Q (new_AGEMA_signal_17315) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_17316) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M21), .Q (new_AGEMA_signal_17317) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_7249), .Q (new_AGEMA_signal_17318) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_17319) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M23), .Q (new_AGEMA_signal_17320) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_7405), .Q (new_AGEMA_signal_17321) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_17322) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M27), .Q (new_AGEMA_signal_17323) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_7409), .Q (new_AGEMA_signal_17324) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_17325) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M24), .Q (new_AGEMA_signal_17326) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_7597), .Q (new_AGEMA_signal_17327) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_7598), .Q (new_AGEMA_signal_17328) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M21), .Q (new_AGEMA_signal_17329) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_7257), .Q (new_AGEMA_signal_17330) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_17331) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M23), .Q (new_AGEMA_signal_17332) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_7413), .Q (new_AGEMA_signal_17333) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_17334) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M27), .Q (new_AGEMA_signal_17335) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_7417), .Q (new_AGEMA_signal_17336) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_17337) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M24), .Q (new_AGEMA_signal_17338) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_17339) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_17340) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M21), .Q (new_AGEMA_signal_17341) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_7265), .Q (new_AGEMA_signal_17342) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_17343) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M23), .Q (new_AGEMA_signal_17344) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_7421), .Q (new_AGEMA_signal_17345) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_17346) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M27), .Q (new_AGEMA_signal_17347) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_7425), .Q (new_AGEMA_signal_17348) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (new_AGEMA_signal_7426), .Q (new_AGEMA_signal_17349) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M24), .Q (new_AGEMA_signal_17350) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_7617), .Q (new_AGEMA_signal_17351) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_7618), .Q (new_AGEMA_signal_17352) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M21), .Q (new_AGEMA_signal_17353) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_7273), .Q (new_AGEMA_signal_17354) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_7274), .Q (new_AGEMA_signal_17355) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M23), .Q (new_AGEMA_signal_17356) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_7429), .Q (new_AGEMA_signal_17357) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_7430), .Q (new_AGEMA_signal_17358) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M27), .Q (new_AGEMA_signal_17359) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_7433), .Q (new_AGEMA_signal_17360) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_7434), .Q (new_AGEMA_signal_17361) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M24), .Q (new_AGEMA_signal_17362) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_7627), .Q (new_AGEMA_signal_17363) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_17364) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_17365) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_7121), .Q (new_AGEMA_signal_17366) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_7122), .Q (new_AGEMA_signal_17367) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_17368) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_7277), .Q (new_AGEMA_signal_17369) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_7278), .Q (new_AGEMA_signal_17370) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_17371) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_7281), .Q (new_AGEMA_signal_17372) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (new_AGEMA_signal_7282), .Q (new_AGEMA_signal_17373) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_17374) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_7437), .Q (new_AGEMA_signal_17375) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_7438), .Q (new_AGEMA_signal_17376) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_17377) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_7129), .Q (new_AGEMA_signal_17378) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_7130), .Q (new_AGEMA_signal_17379) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_17380) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_7285), .Q (new_AGEMA_signal_17381) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_7286), .Q (new_AGEMA_signal_17382) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_17383) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_7289), .Q (new_AGEMA_signal_17384) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_17385) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_17386) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_17387) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_17388) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_17389) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_7137), .Q (new_AGEMA_signal_17390) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_7138), .Q (new_AGEMA_signal_17391) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_17392) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_7293), .Q (new_AGEMA_signal_17393) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_17394) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_17395) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_7297), .Q (new_AGEMA_signal_17396) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_17397) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_17398) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_7457), .Q (new_AGEMA_signal_17399) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_17400) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_17401) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_7145), .Q (new_AGEMA_signal_17402) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_17403) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_17404) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_7301), .Q (new_AGEMA_signal_17405) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_17406) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_17407) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_7305), .Q (new_AGEMA_signal_17408) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_17409) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_17410) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_17411) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_17412) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_17653), .Q (new_AGEMA_signal_17654) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_17657), .Q (new_AGEMA_signal_17658) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_17661), .Q (new_AGEMA_signal_17662) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_17665), .Q (new_AGEMA_signal_17666) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_17669), .Q (new_AGEMA_signal_17670) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_17673), .Q (new_AGEMA_signal_17674) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_17677), .Q (new_AGEMA_signal_17678) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_17681), .Q (new_AGEMA_signal_17682) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_17685), .Q (new_AGEMA_signal_17686) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_17689), .Q (new_AGEMA_signal_17690) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_17693), .Q (new_AGEMA_signal_17694) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_17697), .Q (new_AGEMA_signal_17698) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_17701), .Q (new_AGEMA_signal_17702) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_17705), .Q (new_AGEMA_signal_17706) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_17709), .Q (new_AGEMA_signal_17710) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_17713), .Q (new_AGEMA_signal_17714) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_17717), .Q (new_AGEMA_signal_17718) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_17721), .Q (new_AGEMA_signal_17722) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_17725), .Q (new_AGEMA_signal_17726) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_17729), .Q (new_AGEMA_signal_17730) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_17733), .Q (new_AGEMA_signal_17734) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_17737), .Q (new_AGEMA_signal_17738) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_17741), .Q (new_AGEMA_signal_17742) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_17745), .Q (new_AGEMA_signal_17746) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_17749), .Q (new_AGEMA_signal_17750) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_17753), .Q (new_AGEMA_signal_17754) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_17757), .Q (new_AGEMA_signal_17758) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_17761), .Q (new_AGEMA_signal_17762) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_17765), .Q (new_AGEMA_signal_17766) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_17769), .Q (new_AGEMA_signal_17770) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_17773), .Q (new_AGEMA_signal_17774) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_17777), .Q (new_AGEMA_signal_17778) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_17781), .Q (new_AGEMA_signal_17782) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_17785), .Q (new_AGEMA_signal_17786) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_17789), .Q (new_AGEMA_signal_17790) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_17793), .Q (new_AGEMA_signal_17794) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_17797), .Q (new_AGEMA_signal_17798) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_17801), .Q (new_AGEMA_signal_17802) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_17805), .Q (new_AGEMA_signal_17806) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_17809), .Q (new_AGEMA_signal_17810) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_17813), .Q (new_AGEMA_signal_17814) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_17817), .Q (new_AGEMA_signal_17818) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_17821), .Q (new_AGEMA_signal_17822) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_17825), .Q (new_AGEMA_signal_17826) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_17829), .Q (new_AGEMA_signal_17830) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_17833), .Q (new_AGEMA_signal_17834) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_17837), .Q (new_AGEMA_signal_17838) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_17841), .Q (new_AGEMA_signal_17842) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_17845), .Q (new_AGEMA_signal_17846) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_17849), .Q (new_AGEMA_signal_17850) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_17853), .Q (new_AGEMA_signal_17854) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_17857), .Q (new_AGEMA_signal_17858) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_17861), .Q (new_AGEMA_signal_17862) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_17865), .Q (new_AGEMA_signal_17866) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_17869), .Q (new_AGEMA_signal_17870) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_17873), .Q (new_AGEMA_signal_17874) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_17877), .Q (new_AGEMA_signal_17878) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_17881), .Q (new_AGEMA_signal_17882) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_17885), .Q (new_AGEMA_signal_17886) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_17889), .Q (new_AGEMA_signal_17890) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_17893), .Q (new_AGEMA_signal_17894) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_17897), .Q (new_AGEMA_signal_17898) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_17901), .Q (new_AGEMA_signal_17902) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_17905), .Q (new_AGEMA_signal_17906) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_17909), .Q (new_AGEMA_signal_17910) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_17913), .Q (new_AGEMA_signal_17914) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_17917), .Q (new_AGEMA_signal_17918) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_17921), .Q (new_AGEMA_signal_17922) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_17925), .Q (new_AGEMA_signal_17926) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_17929), .Q (new_AGEMA_signal_17930) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_17933), .Q (new_AGEMA_signal_17934) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_17937), .Q (new_AGEMA_signal_17938) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_17941), .Q (new_AGEMA_signal_17942) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_17945), .Q (new_AGEMA_signal_17946) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_17949), .Q (new_AGEMA_signal_17950) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_17953), .Q (new_AGEMA_signal_17954) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_17957), .Q (new_AGEMA_signal_17958) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_17961), .Q (new_AGEMA_signal_17962) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_17965), .Q (new_AGEMA_signal_17966) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_17969), .Q (new_AGEMA_signal_17970) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_17973), .Q (new_AGEMA_signal_17974) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_17977), .Q (new_AGEMA_signal_17978) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_17981), .Q (new_AGEMA_signal_17982) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_17985), .Q (new_AGEMA_signal_17986) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_17989), .Q (new_AGEMA_signal_17990) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_17993), .Q (new_AGEMA_signal_17994) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_17997), .Q (new_AGEMA_signal_17998) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_18001), .Q (new_AGEMA_signal_18002) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_18005), .Q (new_AGEMA_signal_18006) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_18009), .Q (new_AGEMA_signal_18010) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_18013), .Q (new_AGEMA_signal_18014) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_18017), .Q (new_AGEMA_signal_18018) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_18021), .Q (new_AGEMA_signal_18022) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_18025), .Q (new_AGEMA_signal_18026) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_18029), .Q (new_AGEMA_signal_18030) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_18033), .Q (new_AGEMA_signal_18034) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_18037), .Q (new_AGEMA_signal_18038) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_18041), .Q (new_AGEMA_signal_18042) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_18045), .Q (new_AGEMA_signal_18046) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_18049), .Q (new_AGEMA_signal_18050) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_18053), .Q (new_AGEMA_signal_18054) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_18057), .Q (new_AGEMA_signal_18058) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_18061), .Q (new_AGEMA_signal_18062) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_18065), .Q (new_AGEMA_signal_18066) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_18069), .Q (new_AGEMA_signal_18070) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_18073), .Q (new_AGEMA_signal_18074) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_18077), .Q (new_AGEMA_signal_18078) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_18081), .Q (new_AGEMA_signal_18082) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_18085), .Q (new_AGEMA_signal_18086) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_18089), .Q (new_AGEMA_signal_18090) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_18093), .Q (new_AGEMA_signal_18094) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_18097), .Q (new_AGEMA_signal_18098) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_18101), .Q (new_AGEMA_signal_18102) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_18105), .Q (new_AGEMA_signal_18106) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_18109), .Q (new_AGEMA_signal_18110) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_18113), .Q (new_AGEMA_signal_18114) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_18117), .Q (new_AGEMA_signal_18118) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_18121), .Q (new_AGEMA_signal_18122) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_18125), .Q (new_AGEMA_signal_18126) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_18129), .Q (new_AGEMA_signal_18130) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_18133), .Q (new_AGEMA_signal_18134) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_18137), .Q (new_AGEMA_signal_18138) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_18141), .Q (new_AGEMA_signal_18142) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_18145), .Q (new_AGEMA_signal_18146) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_18149), .Q (new_AGEMA_signal_18150) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_18153), .Q (new_AGEMA_signal_18154) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_18157), .Q (new_AGEMA_signal_18158) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_18161), .Q (new_AGEMA_signal_18162) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_18165), .Q (new_AGEMA_signal_18166) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_18169), .Q (new_AGEMA_signal_18170) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_18173), .Q (new_AGEMA_signal_18174) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_18177), .Q (new_AGEMA_signal_18178) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_18181), .Q (new_AGEMA_signal_18182) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_18185), .Q (new_AGEMA_signal_18186) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_18189), .Q (new_AGEMA_signal_18190) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_18193), .Q (new_AGEMA_signal_18194) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_18197), .Q (new_AGEMA_signal_18198) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_18201), .Q (new_AGEMA_signal_18202) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_18205), .Q (new_AGEMA_signal_18206) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_18209), .Q (new_AGEMA_signal_18210) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_18213), .Q (new_AGEMA_signal_18214) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_18217), .Q (new_AGEMA_signal_18218) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_18221), .Q (new_AGEMA_signal_18222) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_18225), .Q (new_AGEMA_signal_18226) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_18229), .Q (new_AGEMA_signal_18230) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_18233), .Q (new_AGEMA_signal_18234) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_18237), .Q (new_AGEMA_signal_18238) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_18241), .Q (new_AGEMA_signal_18242) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_18245), .Q (new_AGEMA_signal_18246) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_18249), .Q (new_AGEMA_signal_18250) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_18253), .Q (new_AGEMA_signal_18254) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_18257), .Q (new_AGEMA_signal_18258) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_18261), .Q (new_AGEMA_signal_18262) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_18265), .Q (new_AGEMA_signal_18266) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_18269), .Q (new_AGEMA_signal_18270) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_18273), .Q (new_AGEMA_signal_18274) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_18277), .Q (new_AGEMA_signal_18278) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_18281), .Q (new_AGEMA_signal_18282) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_18285), .Q (new_AGEMA_signal_18286) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_18289), .Q (new_AGEMA_signal_18290) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_18293), .Q (new_AGEMA_signal_18294) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_18297), .Q (new_AGEMA_signal_18298) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_18301), .Q (new_AGEMA_signal_18302) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_18305), .Q (new_AGEMA_signal_18306) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_18309), .Q (new_AGEMA_signal_18310) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_18313), .Q (new_AGEMA_signal_18314) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_18317), .Q (new_AGEMA_signal_18318) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_18321), .Q (new_AGEMA_signal_18322) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_18325), .Q (new_AGEMA_signal_18326) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_18329), .Q (new_AGEMA_signal_18330) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_18333), .Q (new_AGEMA_signal_18334) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_18337), .Q (new_AGEMA_signal_18338) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_18341), .Q (new_AGEMA_signal_18342) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_18345), .Q (new_AGEMA_signal_18346) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_18349), .Q (new_AGEMA_signal_18350) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_18353), .Q (new_AGEMA_signal_18354) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_18357), .Q (new_AGEMA_signal_18358) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_18361), .Q (new_AGEMA_signal_18362) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_18365), .Q (new_AGEMA_signal_18366) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_18369), .Q (new_AGEMA_signal_18370) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_18373), .Q (new_AGEMA_signal_18374) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_18377), .Q (new_AGEMA_signal_18378) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_18381), .Q (new_AGEMA_signal_18382) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_18385), .Q (new_AGEMA_signal_18386) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_18389), .Q (new_AGEMA_signal_18390) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_18393), .Q (new_AGEMA_signal_18394) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_18397), .Q (new_AGEMA_signal_18398) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_18401), .Q (new_AGEMA_signal_18402) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_18405), .Q (new_AGEMA_signal_18406) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_18409), .Q (new_AGEMA_signal_18410) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_18413), .Q (new_AGEMA_signal_18414) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_18417), .Q (new_AGEMA_signal_18418) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_18421), .Q (new_AGEMA_signal_18422) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_18425), .Q (new_AGEMA_signal_18426) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_18429), .Q (new_AGEMA_signal_18430) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_18433), .Q (new_AGEMA_signal_18434) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_18437), .Q (new_AGEMA_signal_18438) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_18441), .Q (new_AGEMA_signal_18442) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_18445), .Q (new_AGEMA_signal_18446) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_18449), .Q (new_AGEMA_signal_18450) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_18453), .Q (new_AGEMA_signal_18454) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_18457), .Q (new_AGEMA_signal_18458) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_18461), .Q (new_AGEMA_signal_18462) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_18465), .Q (new_AGEMA_signal_18466) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_18469), .Q (new_AGEMA_signal_18470) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_18473), .Q (new_AGEMA_signal_18474) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_18477), .Q (new_AGEMA_signal_18478) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_18481), .Q (new_AGEMA_signal_18482) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_18485), .Q (new_AGEMA_signal_18486) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_18489), .Q (new_AGEMA_signal_18490) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_18493), .Q (new_AGEMA_signal_18494) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_18497), .Q (new_AGEMA_signal_18498) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_18501), .Q (new_AGEMA_signal_18502) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_18505), .Q (new_AGEMA_signal_18506) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_18509), .Q (new_AGEMA_signal_18510) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_18513), .Q (new_AGEMA_signal_18514) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_18517), .Q (new_AGEMA_signal_18518) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_18521), .Q (new_AGEMA_signal_18522) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_18525), .Q (new_AGEMA_signal_18526) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_18529), .Q (new_AGEMA_signal_18530) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_18533), .Q (new_AGEMA_signal_18534) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_18537), .Q (new_AGEMA_signal_18538) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_18541), .Q (new_AGEMA_signal_18542) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_18545), .Q (new_AGEMA_signal_18546) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_18549), .Q (new_AGEMA_signal_18550) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_18553), .Q (new_AGEMA_signal_18554) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_18557), .Q (new_AGEMA_signal_18558) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_18561), .Q (new_AGEMA_signal_18562) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_18565), .Q (new_AGEMA_signal_18566) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_18569), .Q (new_AGEMA_signal_18570) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_18573), .Q (new_AGEMA_signal_18574) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_18577), .Q (new_AGEMA_signal_18578) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_18581), .Q (new_AGEMA_signal_18582) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_18585), .Q (new_AGEMA_signal_18586) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_18589), .Q (new_AGEMA_signal_18590) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_18593), .Q (new_AGEMA_signal_18594) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_18597), .Q (new_AGEMA_signal_18598) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_18601), .Q (new_AGEMA_signal_18602) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_18605), .Q (new_AGEMA_signal_18606) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_18609), .Q (new_AGEMA_signal_18610) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_18613), .Q (new_AGEMA_signal_18614) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_18617), .Q (new_AGEMA_signal_18618) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_18621), .Q (new_AGEMA_signal_18622) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_18625), .Q (new_AGEMA_signal_18626) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_18629), .Q (new_AGEMA_signal_18630) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_18633), .Q (new_AGEMA_signal_18634) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_18637), .Q (new_AGEMA_signal_18638) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_18641), .Q (new_AGEMA_signal_18642) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_18645), .Q (new_AGEMA_signal_18646) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_18649), .Q (new_AGEMA_signal_18650) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_18653), .Q (new_AGEMA_signal_18654) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_18657), .Q (new_AGEMA_signal_18658) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_18661), .Q (new_AGEMA_signal_18662) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_18665), .Q (new_AGEMA_signal_18666) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_18669), .Q (new_AGEMA_signal_18670) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_18673), .Q (new_AGEMA_signal_18674) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_18677), .Q (new_AGEMA_signal_18678) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_18681), .Q (new_AGEMA_signal_18682) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_18685), .Q (new_AGEMA_signal_18686) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_18689), .Q (new_AGEMA_signal_18690) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_18693), .Q (new_AGEMA_signal_18694) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_18697), .Q (new_AGEMA_signal_18698) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_18701), .Q (new_AGEMA_signal_18702) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_18705), .Q (new_AGEMA_signal_18706) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_18709), .Q (new_AGEMA_signal_18710) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_18713), .Q (new_AGEMA_signal_18714) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_18717), .Q (new_AGEMA_signal_18718) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_18721), .Q (new_AGEMA_signal_18722) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_18725), .Q (new_AGEMA_signal_18726) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_18729), .Q (new_AGEMA_signal_18730) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_18733), .Q (new_AGEMA_signal_18734) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_18737), .Q (new_AGEMA_signal_18738) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_18741), .Q (new_AGEMA_signal_18742) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_18745), .Q (new_AGEMA_signal_18746) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_18749), .Q (new_AGEMA_signal_18750) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_18753), .Q (new_AGEMA_signal_18754) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_18757), .Q (new_AGEMA_signal_18758) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_18761), .Q (new_AGEMA_signal_18762) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_18765), .Q (new_AGEMA_signal_18766) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_18769), .Q (new_AGEMA_signal_18770) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_18773), .Q (new_AGEMA_signal_18774) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_18777), .Q (new_AGEMA_signal_18778) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_18781), .Q (new_AGEMA_signal_18782) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_18785), .Q (new_AGEMA_signal_18786) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_18789), .Q (new_AGEMA_signal_18790) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_18793), .Q (new_AGEMA_signal_18794) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_18797), .Q (new_AGEMA_signal_18798) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_18801), .Q (new_AGEMA_signal_18802) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_18805), .Q (new_AGEMA_signal_18806) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_18809), .Q (new_AGEMA_signal_18810) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_18813), .Q (new_AGEMA_signal_18814) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_18817), .Q (new_AGEMA_signal_18818) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_18821), .Q (new_AGEMA_signal_18822) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_18825), .Q (new_AGEMA_signal_18826) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_18829), .Q (new_AGEMA_signal_18830) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_18833), .Q (new_AGEMA_signal_18834) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_18837), .Q (new_AGEMA_signal_18838) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_18841), .Q (new_AGEMA_signal_18842) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_18845), .Q (new_AGEMA_signal_18846) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_18849), .Q (new_AGEMA_signal_18850) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_18853), .Q (new_AGEMA_signal_18854) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_18857), .Q (new_AGEMA_signal_18858) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_18861), .Q (new_AGEMA_signal_18862) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_18865), .Q (new_AGEMA_signal_18866) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_18869), .Q (new_AGEMA_signal_18870) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_18873), .Q (new_AGEMA_signal_18874) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_18877), .Q (new_AGEMA_signal_18878) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_18881), .Q (new_AGEMA_signal_18882) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_18885), .Q (new_AGEMA_signal_18886) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_18889), .Q (new_AGEMA_signal_18890) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_18893), .Q (new_AGEMA_signal_18894) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_18897), .Q (new_AGEMA_signal_18898) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_18901), .Q (new_AGEMA_signal_18902) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_18905), .Q (new_AGEMA_signal_18906) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_18909), .Q (new_AGEMA_signal_18910) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_18913), .Q (new_AGEMA_signal_18914) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_18917), .Q (new_AGEMA_signal_18918) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_18921), .Q (new_AGEMA_signal_18922) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_18925), .Q (new_AGEMA_signal_18926) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_18929), .Q (new_AGEMA_signal_18930) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_18933), .Q (new_AGEMA_signal_18934) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_18937), .Q (new_AGEMA_signal_18938) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_18941), .Q (new_AGEMA_signal_18942) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_18945), .Q (new_AGEMA_signal_18946) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_18949), .Q (new_AGEMA_signal_18950) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_18953), .Q (new_AGEMA_signal_18954) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_18957), .Q (new_AGEMA_signal_18958) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_18961), .Q (new_AGEMA_signal_18962) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_18965), .Q (new_AGEMA_signal_18966) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_18969), .Q (new_AGEMA_signal_18970) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_18973), .Q (new_AGEMA_signal_18974) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_18977), .Q (new_AGEMA_signal_18978) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_18981), .Q (new_AGEMA_signal_18982) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_18985), .Q (new_AGEMA_signal_18986) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_18989), .Q (new_AGEMA_signal_18990) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_18993), .Q (new_AGEMA_signal_18994) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_18997), .Q (new_AGEMA_signal_18998) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_19001), .Q (new_AGEMA_signal_19002) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_19005), .Q (new_AGEMA_signal_19006) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_19009), .Q (new_AGEMA_signal_19010) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_19013), .Q (new_AGEMA_signal_19014) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_19017), .Q (new_AGEMA_signal_19018) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_19021), .Q (new_AGEMA_signal_19022) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_19025), .Q (new_AGEMA_signal_19026) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_19029), .Q (new_AGEMA_signal_19030) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_19033), .Q (new_AGEMA_signal_19034) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_19037), .Q (new_AGEMA_signal_19038) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_19041), .Q (new_AGEMA_signal_19042) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_19045), .Q (new_AGEMA_signal_19046) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_19049), .Q (new_AGEMA_signal_19050) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_19053), .Q (new_AGEMA_signal_19054) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_19057), .Q (new_AGEMA_signal_19058) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_19061), .Q (new_AGEMA_signal_19062) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_19065), .Q (new_AGEMA_signal_19066) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_19069), .Q (new_AGEMA_signal_19070) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_19073), .Q (new_AGEMA_signal_19074) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_19077), .Q (new_AGEMA_signal_19078) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_19081), .Q (new_AGEMA_signal_19082) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_19085), .Q (new_AGEMA_signal_19086) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_19089), .Q (new_AGEMA_signal_19090) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_19093), .Q (new_AGEMA_signal_19094) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_19097), .Q (new_AGEMA_signal_19098) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_19101), .Q (new_AGEMA_signal_19102) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_19105), .Q (new_AGEMA_signal_19106) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_19109), .Q (new_AGEMA_signal_19110) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_19113), .Q (new_AGEMA_signal_19114) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_19117), .Q (new_AGEMA_signal_19118) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_19121), .Q (new_AGEMA_signal_19122) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_19125), .Q (new_AGEMA_signal_19126) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_19129), .Q (new_AGEMA_signal_19130) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_19133), .Q (new_AGEMA_signal_19134) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_19137), .Q (new_AGEMA_signal_19138) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_19141), .Q (new_AGEMA_signal_19142) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_19145), .Q (new_AGEMA_signal_19146) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_19149), .Q (new_AGEMA_signal_19150) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_19153), .Q (new_AGEMA_signal_19154) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_19157), .Q (new_AGEMA_signal_19158) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_19161), .Q (new_AGEMA_signal_19162) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_19165), .Q (new_AGEMA_signal_19166) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_19169), .Q (new_AGEMA_signal_19170) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_19173), .Q (new_AGEMA_signal_19174) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_19177), .Q (new_AGEMA_signal_19178) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_19181), .Q (new_AGEMA_signal_19182) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_19185), .Q (new_AGEMA_signal_19186) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_19189), .Q (new_AGEMA_signal_19190) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_19193), .Q (new_AGEMA_signal_19194) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_19197), .Q (new_AGEMA_signal_19198) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_19201), .Q (new_AGEMA_signal_19202) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_19205), .Q (new_AGEMA_signal_19206) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_19209), .Q (new_AGEMA_signal_19210) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_19213), .Q (new_AGEMA_signal_19214) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_19217), .Q (new_AGEMA_signal_19218) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_19221), .Q (new_AGEMA_signal_19222) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C (clk), .D (new_AGEMA_signal_19224), .Q (new_AGEMA_signal_19225) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_19227), .Q (new_AGEMA_signal_19228) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C (clk), .D (new_AGEMA_signal_19230), .Q (new_AGEMA_signal_19231) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_19233), .Q (new_AGEMA_signal_19234) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C (clk), .D (new_AGEMA_signal_19236), .Q (new_AGEMA_signal_19237) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C (clk), .D (new_AGEMA_signal_19239), .Q (new_AGEMA_signal_19240) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C (clk), .D (new_AGEMA_signal_19242), .Q (new_AGEMA_signal_19243) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_19245), .Q (new_AGEMA_signal_19246) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C (clk), .D (new_AGEMA_signal_19248), .Q (new_AGEMA_signal_19249) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_19251), .Q (new_AGEMA_signal_19252) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C (clk), .D (new_AGEMA_signal_19254), .Q (new_AGEMA_signal_19255) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_19257), .Q (new_AGEMA_signal_19258) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C (clk), .D (new_AGEMA_signal_19260), .Q (new_AGEMA_signal_19261) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_19263), .Q (new_AGEMA_signal_19264) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C (clk), .D (new_AGEMA_signal_19266), .Q (new_AGEMA_signal_19267) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_19269), .Q (new_AGEMA_signal_19270) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C (clk), .D (new_AGEMA_signal_19272), .Q (new_AGEMA_signal_19273) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_19275), .Q (new_AGEMA_signal_19276) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C (clk), .D (new_AGEMA_signal_19278), .Q (new_AGEMA_signal_19279) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_19281), .Q (new_AGEMA_signal_19282) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C (clk), .D (new_AGEMA_signal_19284), .Q (new_AGEMA_signal_19285) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_19287), .Q (new_AGEMA_signal_19288) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C (clk), .D (new_AGEMA_signal_19290), .Q (new_AGEMA_signal_19291) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_19293), .Q (new_AGEMA_signal_19294) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C (clk), .D (new_AGEMA_signal_19296), .Q (new_AGEMA_signal_19297) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_19299), .Q (new_AGEMA_signal_19300) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C (clk), .D (new_AGEMA_signal_19302), .Q (new_AGEMA_signal_19303) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_19305), .Q (new_AGEMA_signal_19306) ) ;
    buf_clk new_AGEMA_reg_buffer_6585 ( .C (clk), .D (new_AGEMA_signal_19308), .Q (new_AGEMA_signal_19309) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_19311), .Q (new_AGEMA_signal_19312) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C (clk), .D (new_AGEMA_signal_19314), .Q (new_AGEMA_signal_19315) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_19317), .Q (new_AGEMA_signal_19318) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C (clk), .D (new_AGEMA_signal_19320), .Q (new_AGEMA_signal_19321) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_19323), .Q (new_AGEMA_signal_19324) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C (clk), .D (new_AGEMA_signal_19326), .Q (new_AGEMA_signal_19327) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_19329), .Q (new_AGEMA_signal_19330) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C (clk), .D (new_AGEMA_signal_19332), .Q (new_AGEMA_signal_19333) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_19335), .Q (new_AGEMA_signal_19336) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C (clk), .D (new_AGEMA_signal_19338), .Q (new_AGEMA_signal_19339) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_19341), .Q (new_AGEMA_signal_19342) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C (clk), .D (new_AGEMA_signal_19344), .Q (new_AGEMA_signal_19345) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C (clk), .D (new_AGEMA_signal_19347), .Q (new_AGEMA_signal_19348) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C (clk), .D (new_AGEMA_signal_19350), .Q (new_AGEMA_signal_19351) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_19353), .Q (new_AGEMA_signal_19354) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C (clk), .D (new_AGEMA_signal_19356), .Q (new_AGEMA_signal_19357) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_19359), .Q (new_AGEMA_signal_19360) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C (clk), .D (new_AGEMA_signal_19362), .Q (new_AGEMA_signal_19363) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_19365), .Q (new_AGEMA_signal_19366) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C (clk), .D (new_AGEMA_signal_19368), .Q (new_AGEMA_signal_19369) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_19371), .Q (new_AGEMA_signal_19372) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C (clk), .D (new_AGEMA_signal_19374), .Q (new_AGEMA_signal_19375) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_19377), .Q (new_AGEMA_signal_19378) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C (clk), .D (new_AGEMA_signal_19380), .Q (new_AGEMA_signal_19381) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_19383), .Q (new_AGEMA_signal_19384) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C (clk), .D (new_AGEMA_signal_19386), .Q (new_AGEMA_signal_19387) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_19389), .Q (new_AGEMA_signal_19390) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C (clk), .D (new_AGEMA_signal_19392), .Q (new_AGEMA_signal_19393) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_19395), .Q (new_AGEMA_signal_19396) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C (clk), .D (new_AGEMA_signal_19398), .Q (new_AGEMA_signal_19399) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_19401), .Q (new_AGEMA_signal_19402) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C (clk), .D (new_AGEMA_signal_19404), .Q (new_AGEMA_signal_19405) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_19407), .Q (new_AGEMA_signal_19408) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C (clk), .D (new_AGEMA_signal_19410), .Q (new_AGEMA_signal_19411) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C (clk), .D (new_AGEMA_signal_19413), .Q (new_AGEMA_signal_19414) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C (clk), .D (new_AGEMA_signal_19416), .Q (new_AGEMA_signal_19417) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C (clk), .D (new_AGEMA_signal_19419), .Q (new_AGEMA_signal_19420) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C (clk), .D (new_AGEMA_signal_19422), .Q (new_AGEMA_signal_19423) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C (clk), .D (new_AGEMA_signal_19425), .Q (new_AGEMA_signal_19426) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C (clk), .D (new_AGEMA_signal_19428), .Q (new_AGEMA_signal_19429) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C (clk), .D (new_AGEMA_signal_19431), .Q (new_AGEMA_signal_19432) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C (clk), .D (new_AGEMA_signal_19434), .Q (new_AGEMA_signal_19435) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C (clk), .D (new_AGEMA_signal_19437), .Q (new_AGEMA_signal_19438) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C (clk), .D (new_AGEMA_signal_19440), .Q (new_AGEMA_signal_19441) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C (clk), .D (new_AGEMA_signal_19443), .Q (new_AGEMA_signal_19444) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C (clk), .D (new_AGEMA_signal_19446), .Q (new_AGEMA_signal_19447) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C (clk), .D (new_AGEMA_signal_19449), .Q (new_AGEMA_signal_19450) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C (clk), .D (new_AGEMA_signal_19452), .Q (new_AGEMA_signal_19453) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C (clk), .D (new_AGEMA_signal_19455), .Q (new_AGEMA_signal_19456) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C (clk), .D (new_AGEMA_signal_19458), .Q (new_AGEMA_signal_19459) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C (clk), .D (new_AGEMA_signal_19461), .Q (new_AGEMA_signal_19462) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C (clk), .D (new_AGEMA_signal_19464), .Q (new_AGEMA_signal_19465) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C (clk), .D (new_AGEMA_signal_19467), .Q (new_AGEMA_signal_19468) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C (clk), .D (new_AGEMA_signal_19470), .Q (new_AGEMA_signal_19471) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C (clk), .D (new_AGEMA_signal_19473), .Q (new_AGEMA_signal_19474) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C (clk), .D (new_AGEMA_signal_19476), .Q (new_AGEMA_signal_19477) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C (clk), .D (new_AGEMA_signal_19479), .Q (new_AGEMA_signal_19480) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C (clk), .D (new_AGEMA_signal_19482), .Q (new_AGEMA_signal_19483) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C (clk), .D (new_AGEMA_signal_19485), .Q (new_AGEMA_signal_19486) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C (clk), .D (new_AGEMA_signal_19488), .Q (new_AGEMA_signal_19489) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C (clk), .D (new_AGEMA_signal_19491), .Q (new_AGEMA_signal_19492) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C (clk), .D (new_AGEMA_signal_19494), .Q (new_AGEMA_signal_19495) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C (clk), .D (new_AGEMA_signal_19497), .Q (new_AGEMA_signal_19498) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C (clk), .D (new_AGEMA_signal_19500), .Q (new_AGEMA_signal_19501) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C (clk), .D (new_AGEMA_signal_19503), .Q (new_AGEMA_signal_19504) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C (clk), .D (new_AGEMA_signal_19506), .Q (new_AGEMA_signal_19507) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C (clk), .D (new_AGEMA_signal_19509), .Q (new_AGEMA_signal_19510) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C (clk), .D (new_AGEMA_signal_19512), .Q (new_AGEMA_signal_19513) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C (clk), .D (new_AGEMA_signal_19515), .Q (new_AGEMA_signal_19516) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C (clk), .D (new_AGEMA_signal_19518), .Q (new_AGEMA_signal_19519) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C (clk), .D (new_AGEMA_signal_19521), .Q (new_AGEMA_signal_19522) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C (clk), .D (new_AGEMA_signal_19524), .Q (new_AGEMA_signal_19525) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C (clk), .D (new_AGEMA_signal_19527), .Q (new_AGEMA_signal_19528) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C (clk), .D (new_AGEMA_signal_19530), .Q (new_AGEMA_signal_19531) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C (clk), .D (new_AGEMA_signal_19533), .Q (new_AGEMA_signal_19534) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C (clk), .D (new_AGEMA_signal_19536), .Q (new_AGEMA_signal_19537) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C (clk), .D (new_AGEMA_signal_19539), .Q (new_AGEMA_signal_19540) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C (clk), .D (new_AGEMA_signal_19542), .Q (new_AGEMA_signal_19543) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C (clk), .D (new_AGEMA_signal_19545), .Q (new_AGEMA_signal_19546) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C (clk), .D (new_AGEMA_signal_19548), .Q (new_AGEMA_signal_19549) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C (clk), .D (new_AGEMA_signal_19551), .Q (new_AGEMA_signal_19552) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C (clk), .D (new_AGEMA_signal_19554), .Q (new_AGEMA_signal_19555) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C (clk), .D (new_AGEMA_signal_19557), .Q (new_AGEMA_signal_19558) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C (clk), .D (new_AGEMA_signal_19560), .Q (new_AGEMA_signal_19561) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C (clk), .D (new_AGEMA_signal_19563), .Q (new_AGEMA_signal_19564) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C (clk), .D (new_AGEMA_signal_19566), .Q (new_AGEMA_signal_19567) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C (clk), .D (new_AGEMA_signal_19569), .Q (new_AGEMA_signal_19570) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C (clk), .D (new_AGEMA_signal_19572), .Q (new_AGEMA_signal_19573) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C (clk), .D (new_AGEMA_signal_19575), .Q (new_AGEMA_signal_19576) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C (clk), .D (new_AGEMA_signal_19578), .Q (new_AGEMA_signal_19579) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C (clk), .D (new_AGEMA_signal_19581), .Q (new_AGEMA_signal_19582) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C (clk), .D (new_AGEMA_signal_19584), .Q (new_AGEMA_signal_19585) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C (clk), .D (new_AGEMA_signal_19587), .Q (new_AGEMA_signal_19588) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C (clk), .D (new_AGEMA_signal_19590), .Q (new_AGEMA_signal_19591) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C (clk), .D (new_AGEMA_signal_19593), .Q (new_AGEMA_signal_19594) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C (clk), .D (new_AGEMA_signal_19596), .Q (new_AGEMA_signal_19597) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C (clk), .D (new_AGEMA_signal_19599), .Q (new_AGEMA_signal_19600) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C (clk), .D (new_AGEMA_signal_19602), .Q (new_AGEMA_signal_19603) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C (clk), .D (new_AGEMA_signal_19605), .Q (new_AGEMA_signal_19606) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C (clk), .D (new_AGEMA_signal_19608), .Q (new_AGEMA_signal_19609) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C (clk), .D (new_AGEMA_signal_19611), .Q (new_AGEMA_signal_19612) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C (clk), .D (new_AGEMA_signal_19614), .Q (new_AGEMA_signal_19615) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C (clk), .D (new_AGEMA_signal_19617), .Q (new_AGEMA_signal_19618) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C (clk), .D (new_AGEMA_signal_19620), .Q (new_AGEMA_signal_19621) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C (clk), .D (new_AGEMA_signal_19623), .Q (new_AGEMA_signal_19624) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C (clk), .D (new_AGEMA_signal_19626), .Q (new_AGEMA_signal_19627) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C (clk), .D (new_AGEMA_signal_19629), .Q (new_AGEMA_signal_19630) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C (clk), .D (new_AGEMA_signal_19632), .Q (new_AGEMA_signal_19633) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C (clk), .D (new_AGEMA_signal_19635), .Q (new_AGEMA_signal_19636) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C (clk), .D (new_AGEMA_signal_19638), .Q (new_AGEMA_signal_19639) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C (clk), .D (new_AGEMA_signal_19641), .Q (new_AGEMA_signal_19642) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C (clk), .D (new_AGEMA_signal_19644), .Q (new_AGEMA_signal_19645) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C (clk), .D (new_AGEMA_signal_19647), .Q (new_AGEMA_signal_19648) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C (clk), .D (new_AGEMA_signal_19650), .Q (new_AGEMA_signal_19651) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C (clk), .D (new_AGEMA_signal_19653), .Q (new_AGEMA_signal_19654) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C (clk), .D (new_AGEMA_signal_19656), .Q (new_AGEMA_signal_19657) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C (clk), .D (new_AGEMA_signal_19659), .Q (new_AGEMA_signal_19660) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C (clk), .D (new_AGEMA_signal_19662), .Q (new_AGEMA_signal_19663) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C (clk), .D (new_AGEMA_signal_19665), .Q (new_AGEMA_signal_19666) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C (clk), .D (new_AGEMA_signal_19668), .Q (new_AGEMA_signal_19669) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C (clk), .D (new_AGEMA_signal_19671), .Q (new_AGEMA_signal_19672) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C (clk), .D (new_AGEMA_signal_19674), .Q (new_AGEMA_signal_19675) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C (clk), .D (new_AGEMA_signal_19677), .Q (new_AGEMA_signal_19678) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C (clk), .D (new_AGEMA_signal_19680), .Q (new_AGEMA_signal_19681) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C (clk), .D (new_AGEMA_signal_19683), .Q (new_AGEMA_signal_19684) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C (clk), .D (new_AGEMA_signal_19686), .Q (new_AGEMA_signal_19687) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C (clk), .D (new_AGEMA_signal_19689), .Q (new_AGEMA_signal_19690) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C (clk), .D (new_AGEMA_signal_19692), .Q (new_AGEMA_signal_19693) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C (clk), .D (new_AGEMA_signal_19695), .Q (new_AGEMA_signal_19696) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C (clk), .D (new_AGEMA_signal_19698), .Q (new_AGEMA_signal_19699) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C (clk), .D (new_AGEMA_signal_19701), .Q (new_AGEMA_signal_19702) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C (clk), .D (new_AGEMA_signal_19704), .Q (new_AGEMA_signal_19705) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C (clk), .D (new_AGEMA_signal_19707), .Q (new_AGEMA_signal_19708) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C (clk), .D (new_AGEMA_signal_19710), .Q (new_AGEMA_signal_19711) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C (clk), .D (new_AGEMA_signal_19713), .Q (new_AGEMA_signal_19714) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C (clk), .D (new_AGEMA_signal_19716), .Q (new_AGEMA_signal_19717) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C (clk), .D (new_AGEMA_signal_19719), .Q (new_AGEMA_signal_19720) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C (clk), .D (new_AGEMA_signal_19722), .Q (new_AGEMA_signal_19723) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C (clk), .D (new_AGEMA_signal_19725), .Q (new_AGEMA_signal_19726) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C (clk), .D (new_AGEMA_signal_19728), .Q (new_AGEMA_signal_19729) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C (clk), .D (new_AGEMA_signal_19731), .Q (new_AGEMA_signal_19732) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C (clk), .D (new_AGEMA_signal_19734), .Q (new_AGEMA_signal_19735) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C (clk), .D (new_AGEMA_signal_19737), .Q (new_AGEMA_signal_19738) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C (clk), .D (new_AGEMA_signal_19740), .Q (new_AGEMA_signal_19741) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C (clk), .D (new_AGEMA_signal_19743), .Q (new_AGEMA_signal_19744) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C (clk), .D (new_AGEMA_signal_19746), .Q (new_AGEMA_signal_19747) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C (clk), .D (new_AGEMA_signal_19749), .Q (new_AGEMA_signal_19750) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C (clk), .D (new_AGEMA_signal_19752), .Q (new_AGEMA_signal_19753) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C (clk), .D (new_AGEMA_signal_19755), .Q (new_AGEMA_signal_19756) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C (clk), .D (new_AGEMA_signal_19758), .Q (new_AGEMA_signal_19759) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C (clk), .D (new_AGEMA_signal_19761), .Q (new_AGEMA_signal_19762) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C (clk), .D (new_AGEMA_signal_19764), .Q (new_AGEMA_signal_19765) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C (clk), .D (new_AGEMA_signal_19767), .Q (new_AGEMA_signal_19768) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C (clk), .D (new_AGEMA_signal_19770), .Q (new_AGEMA_signal_19771) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C (clk), .D (new_AGEMA_signal_19773), .Q (new_AGEMA_signal_19774) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C (clk), .D (new_AGEMA_signal_19776), .Q (new_AGEMA_signal_19777) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C (clk), .D (new_AGEMA_signal_19779), .Q (new_AGEMA_signal_19780) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C (clk), .D (new_AGEMA_signal_19782), .Q (new_AGEMA_signal_19783) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C (clk), .D (new_AGEMA_signal_19785), .Q (new_AGEMA_signal_19786) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C (clk), .D (new_AGEMA_signal_19788), .Q (new_AGEMA_signal_19789) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C (clk), .D (new_AGEMA_signal_19791), .Q (new_AGEMA_signal_19792) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C (clk), .D (new_AGEMA_signal_19794), .Q (new_AGEMA_signal_19795) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C (clk), .D (new_AGEMA_signal_19797), .Q (new_AGEMA_signal_19798) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C (clk), .D (new_AGEMA_signal_19800), .Q (new_AGEMA_signal_19801) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C (clk), .D (new_AGEMA_signal_19803), .Q (new_AGEMA_signal_19804) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C (clk), .D (new_AGEMA_signal_19806), .Q (new_AGEMA_signal_19807) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C (clk), .D (new_AGEMA_signal_19809), .Q (new_AGEMA_signal_19810) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C (clk), .D (new_AGEMA_signal_19812), .Q (new_AGEMA_signal_19813) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C (clk), .D (new_AGEMA_signal_19815), .Q (new_AGEMA_signal_19816) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C (clk), .D (new_AGEMA_signal_19818), .Q (new_AGEMA_signal_19819) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C (clk), .D (new_AGEMA_signal_19821), .Q (new_AGEMA_signal_19822) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C (clk), .D (new_AGEMA_signal_19824), .Q (new_AGEMA_signal_19825) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C (clk), .D (new_AGEMA_signal_19827), .Q (new_AGEMA_signal_19828) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C (clk), .D (new_AGEMA_signal_19830), .Q (new_AGEMA_signal_19831) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C (clk), .D (new_AGEMA_signal_19833), .Q (new_AGEMA_signal_19834) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C (clk), .D (new_AGEMA_signal_19836), .Q (new_AGEMA_signal_19837) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C (clk), .D (new_AGEMA_signal_19839), .Q (new_AGEMA_signal_19840) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C (clk), .D (new_AGEMA_signal_19842), .Q (new_AGEMA_signal_19843) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C (clk), .D (new_AGEMA_signal_19845), .Q (new_AGEMA_signal_19846) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C (clk), .D (new_AGEMA_signal_19848), .Q (new_AGEMA_signal_19849) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C (clk), .D (new_AGEMA_signal_19851), .Q (new_AGEMA_signal_19852) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C (clk), .D (new_AGEMA_signal_19854), .Q (new_AGEMA_signal_19855) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C (clk), .D (new_AGEMA_signal_19857), .Q (new_AGEMA_signal_19858) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C (clk), .D (new_AGEMA_signal_19860), .Q (new_AGEMA_signal_19861) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C (clk), .D (new_AGEMA_signal_19863), .Q (new_AGEMA_signal_19864) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C (clk), .D (new_AGEMA_signal_19866), .Q (new_AGEMA_signal_19867) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C (clk), .D (new_AGEMA_signal_19869), .Q (new_AGEMA_signal_19870) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C (clk), .D (new_AGEMA_signal_19872), .Q (new_AGEMA_signal_19873) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C (clk), .D (new_AGEMA_signal_19875), .Q (new_AGEMA_signal_19876) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C (clk), .D (new_AGEMA_signal_19878), .Q (new_AGEMA_signal_19879) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C (clk), .D (new_AGEMA_signal_19881), .Q (new_AGEMA_signal_19882) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C (clk), .D (new_AGEMA_signal_19884), .Q (new_AGEMA_signal_19885) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C (clk), .D (new_AGEMA_signal_19887), .Q (new_AGEMA_signal_19888) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C (clk), .D (new_AGEMA_signal_19890), .Q (new_AGEMA_signal_19891) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C (clk), .D (new_AGEMA_signal_19893), .Q (new_AGEMA_signal_19894) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C (clk), .D (new_AGEMA_signal_19896), .Q (new_AGEMA_signal_19897) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C (clk), .D (new_AGEMA_signal_19899), .Q (new_AGEMA_signal_19900) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C (clk), .D (new_AGEMA_signal_19902), .Q (new_AGEMA_signal_19903) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C (clk), .D (new_AGEMA_signal_19905), .Q (new_AGEMA_signal_19906) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C (clk), .D (new_AGEMA_signal_19908), .Q (new_AGEMA_signal_19909) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C (clk), .D (new_AGEMA_signal_19911), .Q (new_AGEMA_signal_19912) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C (clk), .D (new_AGEMA_signal_19914), .Q (new_AGEMA_signal_19915) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C (clk), .D (new_AGEMA_signal_19917), .Q (new_AGEMA_signal_19918) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C (clk), .D (new_AGEMA_signal_19920), .Q (new_AGEMA_signal_19921) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C (clk), .D (new_AGEMA_signal_19923), .Q (new_AGEMA_signal_19924) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C (clk), .D (new_AGEMA_signal_19926), .Q (new_AGEMA_signal_19927) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C (clk), .D (new_AGEMA_signal_19929), .Q (new_AGEMA_signal_19930) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C (clk), .D (new_AGEMA_signal_19932), .Q (new_AGEMA_signal_19933) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C (clk), .D (new_AGEMA_signal_19935), .Q (new_AGEMA_signal_19936) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C (clk), .D (new_AGEMA_signal_19938), .Q (new_AGEMA_signal_19939) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C (clk), .D (new_AGEMA_signal_19941), .Q (new_AGEMA_signal_19942) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C (clk), .D (new_AGEMA_signal_19944), .Q (new_AGEMA_signal_19945) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C (clk), .D (new_AGEMA_signal_19947), .Q (new_AGEMA_signal_19948) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C (clk), .D (new_AGEMA_signal_19950), .Q (new_AGEMA_signal_19951) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C (clk), .D (new_AGEMA_signal_19953), .Q (new_AGEMA_signal_19954) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C (clk), .D (new_AGEMA_signal_19956), .Q (new_AGEMA_signal_19957) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C (clk), .D (new_AGEMA_signal_19959), .Q (new_AGEMA_signal_19960) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C (clk), .D (new_AGEMA_signal_19962), .Q (new_AGEMA_signal_19963) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C (clk), .D (new_AGEMA_signal_19965), .Q (new_AGEMA_signal_19966) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C (clk), .D (new_AGEMA_signal_19968), .Q (new_AGEMA_signal_19969) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C (clk), .D (new_AGEMA_signal_19971), .Q (new_AGEMA_signal_19972) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C (clk), .D (new_AGEMA_signal_19974), .Q (new_AGEMA_signal_19975) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C (clk), .D (new_AGEMA_signal_19977), .Q (new_AGEMA_signal_19978) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C (clk), .D (new_AGEMA_signal_19980), .Q (new_AGEMA_signal_19981) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C (clk), .D (new_AGEMA_signal_19983), .Q (new_AGEMA_signal_19984) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C (clk), .D (new_AGEMA_signal_19986), .Q (new_AGEMA_signal_19987) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C (clk), .D (new_AGEMA_signal_19989), .Q (new_AGEMA_signal_19990) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C (clk), .D (new_AGEMA_signal_19992), .Q (new_AGEMA_signal_19993) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C (clk), .D (new_AGEMA_signal_19995), .Q (new_AGEMA_signal_19996) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C (clk), .D (new_AGEMA_signal_19998), .Q (new_AGEMA_signal_19999) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C (clk), .D (new_AGEMA_signal_20001), .Q (new_AGEMA_signal_20002) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C (clk), .D (new_AGEMA_signal_20004), .Q (new_AGEMA_signal_20005) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C (clk), .D (new_AGEMA_signal_20007), .Q (new_AGEMA_signal_20008) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C (clk), .D (new_AGEMA_signal_20010), .Q (new_AGEMA_signal_20011) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C (clk), .D (new_AGEMA_signal_20013), .Q (new_AGEMA_signal_20014) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C (clk), .D (new_AGEMA_signal_20016), .Q (new_AGEMA_signal_20017) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C (clk), .D (new_AGEMA_signal_20019), .Q (new_AGEMA_signal_20020) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C (clk), .D (new_AGEMA_signal_20022), .Q (new_AGEMA_signal_20023) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C (clk), .D (new_AGEMA_signal_20025), .Q (new_AGEMA_signal_20026) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C (clk), .D (new_AGEMA_signal_20028), .Q (new_AGEMA_signal_20029) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C (clk), .D (new_AGEMA_signal_20031), .Q (new_AGEMA_signal_20032) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C (clk), .D (new_AGEMA_signal_20034), .Q (new_AGEMA_signal_20035) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C (clk), .D (new_AGEMA_signal_20037), .Q (new_AGEMA_signal_20038) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C (clk), .D (new_AGEMA_signal_20040), .Q (new_AGEMA_signal_20041) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C (clk), .D (new_AGEMA_signal_20043), .Q (new_AGEMA_signal_20044) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C (clk), .D (new_AGEMA_signal_20046), .Q (new_AGEMA_signal_20047) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C (clk), .D (new_AGEMA_signal_20049), .Q (new_AGEMA_signal_20050) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C (clk), .D (new_AGEMA_signal_20052), .Q (new_AGEMA_signal_20053) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C (clk), .D (new_AGEMA_signal_20055), .Q (new_AGEMA_signal_20056) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C (clk), .D (new_AGEMA_signal_20058), .Q (new_AGEMA_signal_20059) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C (clk), .D (new_AGEMA_signal_20061), .Q (new_AGEMA_signal_20062) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C (clk), .D (new_AGEMA_signal_20064), .Q (new_AGEMA_signal_20065) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C (clk), .D (new_AGEMA_signal_20067), .Q (new_AGEMA_signal_20068) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C (clk), .D (new_AGEMA_signal_20070), .Q (new_AGEMA_signal_20071) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C (clk), .D (new_AGEMA_signal_20073), .Q (new_AGEMA_signal_20074) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C (clk), .D (new_AGEMA_signal_20076), .Q (new_AGEMA_signal_20077) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C (clk), .D (new_AGEMA_signal_20079), .Q (new_AGEMA_signal_20080) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C (clk), .D (new_AGEMA_signal_20082), .Q (new_AGEMA_signal_20083) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C (clk), .D (new_AGEMA_signal_20085), .Q (new_AGEMA_signal_20086) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C (clk), .D (new_AGEMA_signal_20088), .Q (new_AGEMA_signal_20089) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C (clk), .D (new_AGEMA_signal_20091), .Q (new_AGEMA_signal_20092) ) ;
    buf_clk new_AGEMA_reg_buffer_7371 ( .C (clk), .D (new_AGEMA_signal_20094), .Q (new_AGEMA_signal_20095) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C (clk), .D (new_AGEMA_signal_20097), .Q (new_AGEMA_signal_20098) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C (clk), .D (new_AGEMA_signal_20100), .Q (new_AGEMA_signal_20101) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C (clk), .D (new_AGEMA_signal_20103), .Q (new_AGEMA_signal_20104) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C (clk), .D (new_AGEMA_signal_20106), .Q (new_AGEMA_signal_20107) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C (clk), .D (new_AGEMA_signal_20109), .Q (new_AGEMA_signal_20110) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C (clk), .D (new_AGEMA_signal_20112), .Q (new_AGEMA_signal_20113) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C (clk), .D (new_AGEMA_signal_20115), .Q (new_AGEMA_signal_20116) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C (clk), .D (new_AGEMA_signal_20118), .Q (new_AGEMA_signal_20119) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C (clk), .D (new_AGEMA_signal_20121), .Q (new_AGEMA_signal_20122) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C (clk), .D (new_AGEMA_signal_20124), .Q (new_AGEMA_signal_20125) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C (clk), .D (new_AGEMA_signal_20127), .Q (new_AGEMA_signal_20128) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C (clk), .D (new_AGEMA_signal_20130), .Q (new_AGEMA_signal_20131) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C (clk), .D (new_AGEMA_signal_20133), .Q (new_AGEMA_signal_20134) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C (clk), .D (new_AGEMA_signal_20136), .Q (new_AGEMA_signal_20137) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C (clk), .D (new_AGEMA_signal_20139), .Q (new_AGEMA_signal_20140) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C (clk), .D (new_AGEMA_signal_20142), .Q (new_AGEMA_signal_20143) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C (clk), .D (new_AGEMA_signal_20145), .Q (new_AGEMA_signal_20146) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C (clk), .D (new_AGEMA_signal_20148), .Q (new_AGEMA_signal_20149) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C (clk), .D (new_AGEMA_signal_20151), .Q (new_AGEMA_signal_20152) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C (clk), .D (new_AGEMA_signal_20154), .Q (new_AGEMA_signal_20155) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C (clk), .D (new_AGEMA_signal_20157), .Q (new_AGEMA_signal_20158) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C (clk), .D (new_AGEMA_signal_20160), .Q (new_AGEMA_signal_20161) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C (clk), .D (new_AGEMA_signal_20163), .Q (new_AGEMA_signal_20164) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C (clk), .D (new_AGEMA_signal_20166), .Q (new_AGEMA_signal_20167) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C (clk), .D (new_AGEMA_signal_20169), .Q (new_AGEMA_signal_20170) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C (clk), .D (new_AGEMA_signal_20172), .Q (new_AGEMA_signal_20173) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C (clk), .D (new_AGEMA_signal_20175), .Q (new_AGEMA_signal_20176) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C (clk), .D (new_AGEMA_signal_20178), .Q (new_AGEMA_signal_20179) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C (clk), .D (new_AGEMA_signal_20181), .Q (new_AGEMA_signal_20182) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C (clk), .D (new_AGEMA_signal_20184), .Q (new_AGEMA_signal_20185) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C (clk), .D (new_AGEMA_signal_20187), .Q (new_AGEMA_signal_20188) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C (clk), .D (new_AGEMA_signal_20190), .Q (new_AGEMA_signal_20191) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C (clk), .D (new_AGEMA_signal_20193), .Q (new_AGEMA_signal_20194) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C (clk), .D (new_AGEMA_signal_20196), .Q (new_AGEMA_signal_20197) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C (clk), .D (new_AGEMA_signal_20199), .Q (new_AGEMA_signal_20200) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C (clk), .D (new_AGEMA_signal_20202), .Q (new_AGEMA_signal_20203) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C (clk), .D (new_AGEMA_signal_20205), .Q (new_AGEMA_signal_20206) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C (clk), .D (new_AGEMA_signal_20208), .Q (new_AGEMA_signal_20209) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C (clk), .D (new_AGEMA_signal_20211), .Q (new_AGEMA_signal_20212) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C (clk), .D (new_AGEMA_signal_20214), .Q (new_AGEMA_signal_20215) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C (clk), .D (new_AGEMA_signal_20217), .Q (new_AGEMA_signal_20218) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C (clk), .D (new_AGEMA_signal_20220), .Q (new_AGEMA_signal_20221) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C (clk), .D (new_AGEMA_signal_20223), .Q (new_AGEMA_signal_20224) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C (clk), .D (new_AGEMA_signal_20226), .Q (new_AGEMA_signal_20227) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C (clk), .D (new_AGEMA_signal_20229), .Q (new_AGEMA_signal_20230) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C (clk), .D (new_AGEMA_signal_20232), .Q (new_AGEMA_signal_20233) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C (clk), .D (new_AGEMA_signal_20235), .Q (new_AGEMA_signal_20236) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C (clk), .D (new_AGEMA_signal_20238), .Q (new_AGEMA_signal_20239) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C (clk), .D (new_AGEMA_signal_20241), .Q (new_AGEMA_signal_20242) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C (clk), .D (new_AGEMA_signal_20244), .Q (new_AGEMA_signal_20245) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C (clk), .D (new_AGEMA_signal_20247), .Q (new_AGEMA_signal_20248) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C (clk), .D (new_AGEMA_signal_20250), .Q (new_AGEMA_signal_20251) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C (clk), .D (new_AGEMA_signal_20253), .Q (new_AGEMA_signal_20254) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C (clk), .D (new_AGEMA_signal_20256), .Q (new_AGEMA_signal_20257) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C (clk), .D (new_AGEMA_signal_20259), .Q (new_AGEMA_signal_20260) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C (clk), .D (new_AGEMA_signal_20262), .Q (new_AGEMA_signal_20263) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C (clk), .D (new_AGEMA_signal_20265), .Q (new_AGEMA_signal_20266) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C (clk), .D (new_AGEMA_signal_20268), .Q (new_AGEMA_signal_20269) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C (clk), .D (new_AGEMA_signal_20271), .Q (new_AGEMA_signal_20272) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C (clk), .D (new_AGEMA_signal_20274), .Q (new_AGEMA_signal_20275) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C (clk), .D (new_AGEMA_signal_20277), .Q (new_AGEMA_signal_20278) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C (clk), .D (new_AGEMA_signal_20280), .Q (new_AGEMA_signal_20281) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C (clk), .D (new_AGEMA_signal_20283), .Q (new_AGEMA_signal_20284) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C (clk), .D (new_AGEMA_signal_20286), .Q (new_AGEMA_signal_20287) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C (clk), .D (new_AGEMA_signal_20289), .Q (new_AGEMA_signal_20290) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C (clk), .D (new_AGEMA_signal_20292), .Q (new_AGEMA_signal_20293) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C (clk), .D (new_AGEMA_signal_20295), .Q (new_AGEMA_signal_20296) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C (clk), .D (new_AGEMA_signal_20298), .Q (new_AGEMA_signal_20299) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C (clk), .D (new_AGEMA_signal_20301), .Q (new_AGEMA_signal_20302) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C (clk), .D (new_AGEMA_signal_20304), .Q (new_AGEMA_signal_20305) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C (clk), .D (new_AGEMA_signal_20307), .Q (new_AGEMA_signal_20308) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C (clk), .D (new_AGEMA_signal_20310), .Q (new_AGEMA_signal_20311) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C (clk), .D (new_AGEMA_signal_20313), .Q (new_AGEMA_signal_20314) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C (clk), .D (new_AGEMA_signal_20316), .Q (new_AGEMA_signal_20317) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C (clk), .D (new_AGEMA_signal_20319), .Q (new_AGEMA_signal_20320) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C (clk), .D (new_AGEMA_signal_20322), .Q (new_AGEMA_signal_20323) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C (clk), .D (new_AGEMA_signal_20325), .Q (new_AGEMA_signal_20326) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C (clk), .D (new_AGEMA_signal_20328), .Q (new_AGEMA_signal_20329) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C (clk), .D (new_AGEMA_signal_20331), .Q (new_AGEMA_signal_20332) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C (clk), .D (new_AGEMA_signal_20334), .Q (new_AGEMA_signal_20335) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C (clk), .D (new_AGEMA_signal_20337), .Q (new_AGEMA_signal_20338) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C (clk), .D (new_AGEMA_signal_20340), .Q (new_AGEMA_signal_20341) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C (clk), .D (new_AGEMA_signal_20343), .Q (new_AGEMA_signal_20344) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C (clk), .D (new_AGEMA_signal_20346), .Q (new_AGEMA_signal_20347) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C (clk), .D (new_AGEMA_signal_20349), .Q (new_AGEMA_signal_20350) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C (clk), .D (new_AGEMA_signal_20352), .Q (new_AGEMA_signal_20353) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C (clk), .D (new_AGEMA_signal_20355), .Q (new_AGEMA_signal_20356) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C (clk), .D (new_AGEMA_signal_20358), .Q (new_AGEMA_signal_20359) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C (clk), .D (new_AGEMA_signal_20361), .Q (new_AGEMA_signal_20362) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C (clk), .D (new_AGEMA_signal_20364), .Q (new_AGEMA_signal_20365) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C (clk), .D (new_AGEMA_signal_20367), .Q (new_AGEMA_signal_20368) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C (clk), .D (new_AGEMA_signal_20370), .Q (new_AGEMA_signal_20371) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C (clk), .D (new_AGEMA_signal_20373), .Q (new_AGEMA_signal_20374) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C (clk), .D (new_AGEMA_signal_20376), .Q (new_AGEMA_signal_20377) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C (clk), .D (new_AGEMA_signal_20379), .Q (new_AGEMA_signal_20380) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C (clk), .D (new_AGEMA_signal_20382), .Q (new_AGEMA_signal_20383) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C (clk), .D (new_AGEMA_signal_20385), .Q (new_AGEMA_signal_20386) ) ;
    buf_clk new_AGEMA_reg_buffer_7665 ( .C (clk), .D (new_AGEMA_signal_20388), .Q (new_AGEMA_signal_20389) ) ;
    buf_clk new_AGEMA_reg_buffer_7668 ( .C (clk), .D (new_AGEMA_signal_20391), .Q (new_AGEMA_signal_20392) ) ;
    buf_clk new_AGEMA_reg_buffer_7671 ( .C (clk), .D (new_AGEMA_signal_20394), .Q (new_AGEMA_signal_20395) ) ;
    buf_clk new_AGEMA_reg_buffer_7674 ( .C (clk), .D (new_AGEMA_signal_20397), .Q (new_AGEMA_signal_20398) ) ;
    buf_clk new_AGEMA_reg_buffer_7677 ( .C (clk), .D (new_AGEMA_signal_20400), .Q (new_AGEMA_signal_20401) ) ;
    buf_clk new_AGEMA_reg_buffer_7680 ( .C (clk), .D (new_AGEMA_signal_20403), .Q (new_AGEMA_signal_20404) ) ;
    buf_clk new_AGEMA_reg_buffer_7683 ( .C (clk), .D (new_AGEMA_signal_20406), .Q (new_AGEMA_signal_20407) ) ;
    buf_clk new_AGEMA_reg_buffer_7686 ( .C (clk), .D (new_AGEMA_signal_20409), .Q (new_AGEMA_signal_20410) ) ;
    buf_clk new_AGEMA_reg_buffer_7689 ( .C (clk), .D (new_AGEMA_signal_20412), .Q (new_AGEMA_signal_20413) ) ;
    buf_clk new_AGEMA_reg_buffer_7692 ( .C (clk), .D (new_AGEMA_signal_20415), .Q (new_AGEMA_signal_20416) ) ;
    buf_clk new_AGEMA_reg_buffer_7695 ( .C (clk), .D (new_AGEMA_signal_20418), .Q (new_AGEMA_signal_20419) ) ;
    buf_clk new_AGEMA_reg_buffer_7698 ( .C (clk), .D (new_AGEMA_signal_20421), .Q (new_AGEMA_signal_20422) ) ;
    buf_clk new_AGEMA_reg_buffer_7701 ( .C (clk), .D (new_AGEMA_signal_20424), .Q (new_AGEMA_signal_20425) ) ;
    buf_clk new_AGEMA_reg_buffer_7704 ( .C (clk), .D (new_AGEMA_signal_20427), .Q (new_AGEMA_signal_20428) ) ;
    buf_clk new_AGEMA_reg_buffer_7707 ( .C (clk), .D (new_AGEMA_signal_20430), .Q (new_AGEMA_signal_20431) ) ;
    buf_clk new_AGEMA_reg_buffer_7710 ( .C (clk), .D (new_AGEMA_signal_20433), .Q (new_AGEMA_signal_20434) ) ;
    buf_clk new_AGEMA_reg_buffer_7713 ( .C (clk), .D (new_AGEMA_signal_20436), .Q (new_AGEMA_signal_20437) ) ;
    buf_clk new_AGEMA_reg_buffer_7716 ( .C (clk), .D (new_AGEMA_signal_20439), .Q (new_AGEMA_signal_20440) ) ;
    buf_clk new_AGEMA_reg_buffer_7719 ( .C (clk), .D (new_AGEMA_signal_20442), .Q (new_AGEMA_signal_20443) ) ;
    buf_clk new_AGEMA_reg_buffer_7722 ( .C (clk), .D (new_AGEMA_signal_20445), .Q (new_AGEMA_signal_20446) ) ;
    buf_clk new_AGEMA_reg_buffer_7725 ( .C (clk), .D (new_AGEMA_signal_20448), .Q (new_AGEMA_signal_20449) ) ;
    buf_clk new_AGEMA_reg_buffer_7728 ( .C (clk), .D (new_AGEMA_signal_20451), .Q (new_AGEMA_signal_20452) ) ;
    buf_clk new_AGEMA_reg_buffer_7731 ( .C (clk), .D (new_AGEMA_signal_20454), .Q (new_AGEMA_signal_20455) ) ;
    buf_clk new_AGEMA_reg_buffer_7734 ( .C (clk), .D (new_AGEMA_signal_20457), .Q (new_AGEMA_signal_20458) ) ;
    buf_clk new_AGEMA_reg_buffer_7737 ( .C (clk), .D (new_AGEMA_signal_20460), .Q (new_AGEMA_signal_20461) ) ;
    buf_clk new_AGEMA_reg_buffer_7740 ( .C (clk), .D (new_AGEMA_signal_20463), .Q (new_AGEMA_signal_20464) ) ;
    buf_clk new_AGEMA_reg_buffer_7743 ( .C (clk), .D (new_AGEMA_signal_20466), .Q (new_AGEMA_signal_20467) ) ;
    buf_clk new_AGEMA_reg_buffer_7746 ( .C (clk), .D (new_AGEMA_signal_20469), .Q (new_AGEMA_signal_20470) ) ;
    buf_clk new_AGEMA_reg_buffer_7749 ( .C (clk), .D (new_AGEMA_signal_20472), .Q (new_AGEMA_signal_20473) ) ;
    buf_clk new_AGEMA_reg_buffer_7752 ( .C (clk), .D (new_AGEMA_signal_20475), .Q (new_AGEMA_signal_20476) ) ;
    buf_clk new_AGEMA_reg_buffer_7755 ( .C (clk), .D (new_AGEMA_signal_20478), .Q (new_AGEMA_signal_20479) ) ;
    buf_clk new_AGEMA_reg_buffer_7758 ( .C (clk), .D (new_AGEMA_signal_20481), .Q (new_AGEMA_signal_20482) ) ;
    buf_clk new_AGEMA_reg_buffer_7761 ( .C (clk), .D (new_AGEMA_signal_20484), .Q (new_AGEMA_signal_20485) ) ;
    buf_clk new_AGEMA_reg_buffer_7764 ( .C (clk), .D (new_AGEMA_signal_20487), .Q (new_AGEMA_signal_20488) ) ;
    buf_clk new_AGEMA_reg_buffer_7767 ( .C (clk), .D (new_AGEMA_signal_20490), .Q (new_AGEMA_signal_20491) ) ;
    buf_clk new_AGEMA_reg_buffer_7770 ( .C (clk), .D (new_AGEMA_signal_20493), .Q (new_AGEMA_signal_20494) ) ;
    buf_clk new_AGEMA_reg_buffer_7773 ( .C (clk), .D (new_AGEMA_signal_20496), .Q (new_AGEMA_signal_20497) ) ;
    buf_clk new_AGEMA_reg_buffer_7776 ( .C (clk), .D (new_AGEMA_signal_20499), .Q (new_AGEMA_signal_20500) ) ;
    buf_clk new_AGEMA_reg_buffer_7779 ( .C (clk), .D (new_AGEMA_signal_20502), .Q (new_AGEMA_signal_20503) ) ;
    buf_clk new_AGEMA_reg_buffer_7782 ( .C (clk), .D (new_AGEMA_signal_20505), .Q (new_AGEMA_signal_20506) ) ;
    buf_clk new_AGEMA_reg_buffer_7785 ( .C (clk), .D (new_AGEMA_signal_20508), .Q (new_AGEMA_signal_20509) ) ;
    buf_clk new_AGEMA_reg_buffer_7788 ( .C (clk), .D (new_AGEMA_signal_20511), .Q (new_AGEMA_signal_20512) ) ;
    buf_clk new_AGEMA_reg_buffer_7791 ( .C (clk), .D (new_AGEMA_signal_20514), .Q (new_AGEMA_signal_20515) ) ;
    buf_clk new_AGEMA_reg_buffer_7794 ( .C (clk), .D (new_AGEMA_signal_20517), .Q (new_AGEMA_signal_20518) ) ;
    buf_clk new_AGEMA_reg_buffer_7797 ( .C (clk), .D (new_AGEMA_signal_20520), .Q (new_AGEMA_signal_20521) ) ;
    buf_clk new_AGEMA_reg_buffer_7800 ( .C (clk), .D (new_AGEMA_signal_20523), .Q (new_AGEMA_signal_20524) ) ;
    buf_clk new_AGEMA_reg_buffer_7803 ( .C (clk), .D (new_AGEMA_signal_20526), .Q (new_AGEMA_signal_20527) ) ;
    buf_clk new_AGEMA_reg_buffer_7806 ( .C (clk), .D (new_AGEMA_signal_20529), .Q (new_AGEMA_signal_20530) ) ;
    buf_clk new_AGEMA_reg_buffer_7809 ( .C (clk), .D (new_AGEMA_signal_20532), .Q (new_AGEMA_signal_20533) ) ;
    buf_clk new_AGEMA_reg_buffer_7812 ( .C (clk), .D (new_AGEMA_signal_20535), .Q (new_AGEMA_signal_20536) ) ;
    buf_clk new_AGEMA_reg_buffer_7815 ( .C (clk), .D (new_AGEMA_signal_20538), .Q (new_AGEMA_signal_20539) ) ;
    buf_clk new_AGEMA_reg_buffer_7818 ( .C (clk), .D (new_AGEMA_signal_20541), .Q (new_AGEMA_signal_20542) ) ;
    buf_clk new_AGEMA_reg_buffer_7821 ( .C (clk), .D (new_AGEMA_signal_20544), .Q (new_AGEMA_signal_20545) ) ;
    buf_clk new_AGEMA_reg_buffer_7824 ( .C (clk), .D (new_AGEMA_signal_20547), .Q (new_AGEMA_signal_20548) ) ;
    buf_clk new_AGEMA_reg_buffer_7827 ( .C (clk), .D (new_AGEMA_signal_20550), .Q (new_AGEMA_signal_20551) ) ;
    buf_clk new_AGEMA_reg_buffer_7830 ( .C (clk), .D (new_AGEMA_signal_20553), .Q (new_AGEMA_signal_20554) ) ;
    buf_clk new_AGEMA_reg_buffer_7833 ( .C (clk), .D (new_AGEMA_signal_20556), .Q (new_AGEMA_signal_20557) ) ;
    buf_clk new_AGEMA_reg_buffer_7836 ( .C (clk), .D (new_AGEMA_signal_20559), .Q (new_AGEMA_signal_20560) ) ;
    buf_clk new_AGEMA_reg_buffer_7839 ( .C (clk), .D (new_AGEMA_signal_20562), .Q (new_AGEMA_signal_20563) ) ;
    buf_clk new_AGEMA_reg_buffer_7842 ( .C (clk), .D (new_AGEMA_signal_20565), .Q (new_AGEMA_signal_20566) ) ;
    buf_clk new_AGEMA_reg_buffer_7845 ( .C (clk), .D (new_AGEMA_signal_20568), .Q (new_AGEMA_signal_20569) ) ;
    buf_clk new_AGEMA_reg_buffer_7848 ( .C (clk), .D (new_AGEMA_signal_20571), .Q (new_AGEMA_signal_20572) ) ;
    buf_clk new_AGEMA_reg_buffer_7851 ( .C (clk), .D (new_AGEMA_signal_20574), .Q (new_AGEMA_signal_20575) ) ;
    buf_clk new_AGEMA_reg_buffer_7854 ( .C (clk), .D (new_AGEMA_signal_20577), .Q (new_AGEMA_signal_20578) ) ;
    buf_clk new_AGEMA_reg_buffer_7857 ( .C (clk), .D (new_AGEMA_signal_20580), .Q (new_AGEMA_signal_20581) ) ;
    buf_clk new_AGEMA_reg_buffer_7860 ( .C (clk), .D (new_AGEMA_signal_20583), .Q (new_AGEMA_signal_20584) ) ;
    buf_clk new_AGEMA_reg_buffer_7863 ( .C (clk), .D (new_AGEMA_signal_20586), .Q (new_AGEMA_signal_20587) ) ;
    buf_clk new_AGEMA_reg_buffer_7866 ( .C (clk), .D (new_AGEMA_signal_20589), .Q (new_AGEMA_signal_20590) ) ;
    buf_clk new_AGEMA_reg_buffer_7869 ( .C (clk), .D (new_AGEMA_signal_20592), .Q (new_AGEMA_signal_20593) ) ;
    buf_clk new_AGEMA_reg_buffer_7872 ( .C (clk), .D (new_AGEMA_signal_20595), .Q (new_AGEMA_signal_20596) ) ;
    buf_clk new_AGEMA_reg_buffer_7875 ( .C (clk), .D (new_AGEMA_signal_20598), .Q (new_AGEMA_signal_20599) ) ;
    buf_clk new_AGEMA_reg_buffer_7878 ( .C (clk), .D (new_AGEMA_signal_20601), .Q (new_AGEMA_signal_20602) ) ;
    buf_clk new_AGEMA_reg_buffer_7881 ( .C (clk), .D (new_AGEMA_signal_20604), .Q (new_AGEMA_signal_20605) ) ;
    buf_clk new_AGEMA_reg_buffer_7884 ( .C (clk), .D (new_AGEMA_signal_20607), .Q (new_AGEMA_signal_20608) ) ;
    buf_clk new_AGEMA_reg_buffer_7887 ( .C (clk), .D (new_AGEMA_signal_20610), .Q (new_AGEMA_signal_20611) ) ;
    buf_clk new_AGEMA_reg_buffer_7890 ( .C (clk), .D (new_AGEMA_signal_20613), .Q (new_AGEMA_signal_20614) ) ;
    buf_clk new_AGEMA_reg_buffer_7893 ( .C (clk), .D (new_AGEMA_signal_20616), .Q (new_AGEMA_signal_20617) ) ;
    buf_clk new_AGEMA_reg_buffer_7896 ( .C (clk), .D (new_AGEMA_signal_20619), .Q (new_AGEMA_signal_20620) ) ;
    buf_clk new_AGEMA_reg_buffer_7899 ( .C (clk), .D (new_AGEMA_signal_20622), .Q (new_AGEMA_signal_20623) ) ;
    buf_clk new_AGEMA_reg_buffer_7902 ( .C (clk), .D (new_AGEMA_signal_20625), .Q (new_AGEMA_signal_20626) ) ;
    buf_clk new_AGEMA_reg_buffer_7905 ( .C (clk), .D (new_AGEMA_signal_20628), .Q (new_AGEMA_signal_20629) ) ;
    buf_clk new_AGEMA_reg_buffer_7908 ( .C (clk), .D (new_AGEMA_signal_20631), .Q (new_AGEMA_signal_20632) ) ;
    buf_clk new_AGEMA_reg_buffer_7911 ( .C (clk), .D (new_AGEMA_signal_20634), .Q (new_AGEMA_signal_20635) ) ;
    buf_clk new_AGEMA_reg_buffer_7914 ( .C (clk), .D (new_AGEMA_signal_20637), .Q (new_AGEMA_signal_20638) ) ;
    buf_clk new_AGEMA_reg_buffer_7917 ( .C (clk), .D (new_AGEMA_signal_20640), .Q (new_AGEMA_signal_20641) ) ;
    buf_clk new_AGEMA_reg_buffer_7920 ( .C (clk), .D (new_AGEMA_signal_20643), .Q (new_AGEMA_signal_20644) ) ;
    buf_clk new_AGEMA_reg_buffer_7923 ( .C (clk), .D (new_AGEMA_signal_20646), .Q (new_AGEMA_signal_20647) ) ;
    buf_clk new_AGEMA_reg_buffer_7926 ( .C (clk), .D (new_AGEMA_signal_20649), .Q (new_AGEMA_signal_20650) ) ;
    buf_clk new_AGEMA_reg_buffer_7929 ( .C (clk), .D (new_AGEMA_signal_20652), .Q (new_AGEMA_signal_20653) ) ;
    buf_clk new_AGEMA_reg_buffer_7932 ( .C (clk), .D (new_AGEMA_signal_20655), .Q (new_AGEMA_signal_20656) ) ;
    buf_clk new_AGEMA_reg_buffer_7935 ( .C (clk), .D (new_AGEMA_signal_20658), .Q (new_AGEMA_signal_20659) ) ;
    buf_clk new_AGEMA_reg_buffer_7938 ( .C (clk), .D (new_AGEMA_signal_20661), .Q (new_AGEMA_signal_20662) ) ;
    buf_clk new_AGEMA_reg_buffer_7941 ( .C (clk), .D (new_AGEMA_signal_20664), .Q (new_AGEMA_signal_20665) ) ;
    buf_clk new_AGEMA_reg_buffer_7944 ( .C (clk), .D (new_AGEMA_signal_20667), .Q (new_AGEMA_signal_20668) ) ;
    buf_clk new_AGEMA_reg_buffer_7947 ( .C (clk), .D (new_AGEMA_signal_20670), .Q (new_AGEMA_signal_20671) ) ;
    buf_clk new_AGEMA_reg_buffer_7950 ( .C (clk), .D (new_AGEMA_signal_20673), .Q (new_AGEMA_signal_20674) ) ;
    buf_clk new_AGEMA_reg_buffer_7953 ( .C (clk), .D (new_AGEMA_signal_20676), .Q (new_AGEMA_signal_20677) ) ;
    buf_clk new_AGEMA_reg_buffer_7956 ( .C (clk), .D (new_AGEMA_signal_20679), .Q (new_AGEMA_signal_20680) ) ;
    buf_clk new_AGEMA_reg_buffer_7959 ( .C (clk), .D (new_AGEMA_signal_20682), .Q (new_AGEMA_signal_20683) ) ;
    buf_clk new_AGEMA_reg_buffer_7962 ( .C (clk), .D (new_AGEMA_signal_20685), .Q (new_AGEMA_signal_20686) ) ;
    buf_clk new_AGEMA_reg_buffer_7965 ( .C (clk), .D (new_AGEMA_signal_20688), .Q (new_AGEMA_signal_20689) ) ;
    buf_clk new_AGEMA_reg_buffer_7968 ( .C (clk), .D (new_AGEMA_signal_20691), .Q (new_AGEMA_signal_20692) ) ;
    buf_clk new_AGEMA_reg_buffer_7971 ( .C (clk), .D (new_AGEMA_signal_20694), .Q (new_AGEMA_signal_20695) ) ;
    buf_clk new_AGEMA_reg_buffer_7974 ( .C (clk), .D (new_AGEMA_signal_20697), .Q (new_AGEMA_signal_20698) ) ;
    buf_clk new_AGEMA_reg_buffer_7977 ( .C (clk), .D (new_AGEMA_signal_20700), .Q (new_AGEMA_signal_20701) ) ;
    buf_clk new_AGEMA_reg_buffer_7980 ( .C (clk), .D (new_AGEMA_signal_20703), .Q (new_AGEMA_signal_20704) ) ;
    buf_clk new_AGEMA_reg_buffer_7983 ( .C (clk), .D (new_AGEMA_signal_20706), .Q (new_AGEMA_signal_20707) ) ;
    buf_clk new_AGEMA_reg_buffer_7986 ( .C (clk), .D (new_AGEMA_signal_20709), .Q (new_AGEMA_signal_20710) ) ;
    buf_clk new_AGEMA_reg_buffer_7989 ( .C (clk), .D (new_AGEMA_signal_20712), .Q (new_AGEMA_signal_20713) ) ;
    buf_clk new_AGEMA_reg_buffer_7992 ( .C (clk), .D (new_AGEMA_signal_20715), .Q (new_AGEMA_signal_20716) ) ;
    buf_clk new_AGEMA_reg_buffer_7995 ( .C (clk), .D (new_AGEMA_signal_20718), .Q (new_AGEMA_signal_20719) ) ;
    buf_clk new_AGEMA_reg_buffer_7998 ( .C (clk), .D (new_AGEMA_signal_20721), .Q (new_AGEMA_signal_20722) ) ;
    buf_clk new_AGEMA_reg_buffer_8001 ( .C (clk), .D (new_AGEMA_signal_20724), .Q (new_AGEMA_signal_20725) ) ;
    buf_clk new_AGEMA_reg_buffer_8004 ( .C (clk), .D (new_AGEMA_signal_20727), .Q (new_AGEMA_signal_20728) ) ;
    buf_clk new_AGEMA_reg_buffer_8007 ( .C (clk), .D (new_AGEMA_signal_20730), .Q (new_AGEMA_signal_20731) ) ;
    buf_clk new_AGEMA_reg_buffer_8010 ( .C (clk), .D (new_AGEMA_signal_20733), .Q (new_AGEMA_signal_20734) ) ;
    buf_clk new_AGEMA_reg_buffer_8013 ( .C (clk), .D (new_AGEMA_signal_20736), .Q (new_AGEMA_signal_20737) ) ;
    buf_clk new_AGEMA_reg_buffer_8016 ( .C (clk), .D (new_AGEMA_signal_20739), .Q (new_AGEMA_signal_20740) ) ;
    buf_clk new_AGEMA_reg_buffer_8019 ( .C (clk), .D (new_AGEMA_signal_20742), .Q (new_AGEMA_signal_20743) ) ;
    buf_clk new_AGEMA_reg_buffer_8022 ( .C (clk), .D (new_AGEMA_signal_20745), .Q (new_AGEMA_signal_20746) ) ;
    buf_clk new_AGEMA_reg_buffer_8025 ( .C (clk), .D (new_AGEMA_signal_20748), .Q (new_AGEMA_signal_20749) ) ;
    buf_clk new_AGEMA_reg_buffer_8028 ( .C (clk), .D (new_AGEMA_signal_20751), .Q (new_AGEMA_signal_20752) ) ;
    buf_clk new_AGEMA_reg_buffer_8031 ( .C (clk), .D (new_AGEMA_signal_20754), .Q (new_AGEMA_signal_20755) ) ;
    buf_clk new_AGEMA_reg_buffer_8034 ( .C (clk), .D (new_AGEMA_signal_20757), .Q (new_AGEMA_signal_20758) ) ;
    buf_clk new_AGEMA_reg_buffer_8037 ( .C (clk), .D (new_AGEMA_signal_20760), .Q (new_AGEMA_signal_20761) ) ;
    buf_clk new_AGEMA_reg_buffer_8040 ( .C (clk), .D (new_AGEMA_signal_20763), .Q (new_AGEMA_signal_20764) ) ;
    buf_clk new_AGEMA_reg_buffer_8043 ( .C (clk), .D (new_AGEMA_signal_20766), .Q (new_AGEMA_signal_20767) ) ;
    buf_clk new_AGEMA_reg_buffer_8046 ( .C (clk), .D (new_AGEMA_signal_20769), .Q (new_AGEMA_signal_20770) ) ;
    buf_clk new_AGEMA_reg_buffer_8049 ( .C (clk), .D (new_AGEMA_signal_20772), .Q (new_AGEMA_signal_20773) ) ;
    buf_clk new_AGEMA_reg_buffer_8052 ( .C (clk), .D (new_AGEMA_signal_20775), .Q (new_AGEMA_signal_20776) ) ;
    buf_clk new_AGEMA_reg_buffer_8055 ( .C (clk), .D (new_AGEMA_signal_20778), .Q (new_AGEMA_signal_20779) ) ;
    buf_clk new_AGEMA_reg_buffer_8058 ( .C (clk), .D (new_AGEMA_signal_20781), .Q (new_AGEMA_signal_20782) ) ;
    buf_clk new_AGEMA_reg_buffer_8061 ( .C (clk), .D (new_AGEMA_signal_20784), .Q (new_AGEMA_signal_20785) ) ;
    buf_clk new_AGEMA_reg_buffer_8064 ( .C (clk), .D (new_AGEMA_signal_20787), .Q (new_AGEMA_signal_20788) ) ;
    buf_clk new_AGEMA_reg_buffer_8067 ( .C (clk), .D (new_AGEMA_signal_20790), .Q (new_AGEMA_signal_20791) ) ;
    buf_clk new_AGEMA_reg_buffer_8070 ( .C (clk), .D (new_AGEMA_signal_20793), .Q (new_AGEMA_signal_20794) ) ;
    buf_clk new_AGEMA_reg_buffer_8073 ( .C (clk), .D (new_AGEMA_signal_20796), .Q (new_AGEMA_signal_20797) ) ;
    buf_clk new_AGEMA_reg_buffer_8076 ( .C (clk), .D (new_AGEMA_signal_20799), .Q (new_AGEMA_signal_20800) ) ;
    buf_clk new_AGEMA_reg_buffer_8079 ( .C (clk), .D (new_AGEMA_signal_20802), .Q (new_AGEMA_signal_20803) ) ;
    buf_clk new_AGEMA_reg_buffer_8082 ( .C (clk), .D (new_AGEMA_signal_20805), .Q (new_AGEMA_signal_20806) ) ;
    buf_clk new_AGEMA_reg_buffer_8085 ( .C (clk), .D (new_AGEMA_signal_20808), .Q (new_AGEMA_signal_20809) ) ;
    buf_clk new_AGEMA_reg_buffer_8088 ( .C (clk), .D (new_AGEMA_signal_20811), .Q (new_AGEMA_signal_20812) ) ;
    buf_clk new_AGEMA_reg_buffer_8091 ( .C (clk), .D (new_AGEMA_signal_20814), .Q (new_AGEMA_signal_20815) ) ;
    buf_clk new_AGEMA_reg_buffer_8094 ( .C (clk), .D (new_AGEMA_signal_20817), .Q (new_AGEMA_signal_20818) ) ;
    buf_clk new_AGEMA_reg_buffer_8097 ( .C (clk), .D (new_AGEMA_signal_20820), .Q (new_AGEMA_signal_20821) ) ;
    buf_clk new_AGEMA_reg_buffer_8100 ( .C (clk), .D (new_AGEMA_signal_20823), .Q (new_AGEMA_signal_20824) ) ;
    buf_clk new_AGEMA_reg_buffer_8103 ( .C (clk), .D (new_AGEMA_signal_20826), .Q (new_AGEMA_signal_20827) ) ;
    buf_clk new_AGEMA_reg_buffer_8106 ( .C (clk), .D (new_AGEMA_signal_20829), .Q (new_AGEMA_signal_20830) ) ;
    buf_clk new_AGEMA_reg_buffer_8109 ( .C (clk), .D (new_AGEMA_signal_20832), .Q (new_AGEMA_signal_20833) ) ;
    buf_clk new_AGEMA_reg_buffer_8112 ( .C (clk), .D (new_AGEMA_signal_20835), .Q (new_AGEMA_signal_20836) ) ;
    buf_clk new_AGEMA_reg_buffer_8115 ( .C (clk), .D (new_AGEMA_signal_20838), .Q (new_AGEMA_signal_20839) ) ;
    buf_clk new_AGEMA_reg_buffer_8118 ( .C (clk), .D (new_AGEMA_signal_20841), .Q (new_AGEMA_signal_20842) ) ;
    buf_clk new_AGEMA_reg_buffer_8121 ( .C (clk), .D (new_AGEMA_signal_20844), .Q (new_AGEMA_signal_20845) ) ;
    buf_clk new_AGEMA_reg_buffer_8124 ( .C (clk), .D (new_AGEMA_signal_20847), .Q (new_AGEMA_signal_20848) ) ;
    buf_clk new_AGEMA_reg_buffer_8127 ( .C (clk), .D (new_AGEMA_signal_20850), .Q (new_AGEMA_signal_20851) ) ;
    buf_clk new_AGEMA_reg_buffer_8130 ( .C (clk), .D (new_AGEMA_signal_20853), .Q (new_AGEMA_signal_20854) ) ;
    buf_clk new_AGEMA_reg_buffer_8133 ( .C (clk), .D (new_AGEMA_signal_20856), .Q (new_AGEMA_signal_20857) ) ;
    buf_clk new_AGEMA_reg_buffer_8136 ( .C (clk), .D (new_AGEMA_signal_20859), .Q (new_AGEMA_signal_20860) ) ;
    buf_clk new_AGEMA_reg_buffer_8139 ( .C (clk), .D (new_AGEMA_signal_20862), .Q (new_AGEMA_signal_20863) ) ;
    buf_clk new_AGEMA_reg_buffer_8142 ( .C (clk), .D (new_AGEMA_signal_20865), .Q (new_AGEMA_signal_20866) ) ;
    buf_clk new_AGEMA_reg_buffer_8145 ( .C (clk), .D (new_AGEMA_signal_20868), .Q (new_AGEMA_signal_20869) ) ;
    buf_clk new_AGEMA_reg_buffer_8148 ( .C (clk), .D (new_AGEMA_signal_20871), .Q (new_AGEMA_signal_20872) ) ;
    buf_clk new_AGEMA_reg_buffer_8151 ( .C (clk), .D (new_AGEMA_signal_20874), .Q (new_AGEMA_signal_20875) ) ;
    buf_clk new_AGEMA_reg_buffer_8154 ( .C (clk), .D (new_AGEMA_signal_20877), .Q (new_AGEMA_signal_20878) ) ;
    buf_clk new_AGEMA_reg_buffer_8157 ( .C (clk), .D (new_AGEMA_signal_20880), .Q (new_AGEMA_signal_20881) ) ;
    buf_clk new_AGEMA_reg_buffer_8160 ( .C (clk), .D (new_AGEMA_signal_20883), .Q (new_AGEMA_signal_20884) ) ;
    buf_clk new_AGEMA_reg_buffer_8163 ( .C (clk), .D (new_AGEMA_signal_20886), .Q (new_AGEMA_signal_20887) ) ;
    buf_clk new_AGEMA_reg_buffer_8166 ( .C (clk), .D (new_AGEMA_signal_20889), .Q (new_AGEMA_signal_20890) ) ;
    buf_clk new_AGEMA_reg_buffer_8169 ( .C (clk), .D (new_AGEMA_signal_20892), .Q (new_AGEMA_signal_20893) ) ;
    buf_clk new_AGEMA_reg_buffer_8172 ( .C (clk), .D (new_AGEMA_signal_20895), .Q (new_AGEMA_signal_20896) ) ;
    buf_clk new_AGEMA_reg_buffer_8175 ( .C (clk), .D (new_AGEMA_signal_20898), .Q (new_AGEMA_signal_20899) ) ;
    buf_clk new_AGEMA_reg_buffer_8178 ( .C (clk), .D (new_AGEMA_signal_20901), .Q (new_AGEMA_signal_20902) ) ;
    buf_clk new_AGEMA_reg_buffer_8181 ( .C (clk), .D (new_AGEMA_signal_20904), .Q (new_AGEMA_signal_20905) ) ;
    buf_clk new_AGEMA_reg_buffer_8184 ( .C (clk), .D (new_AGEMA_signal_20907), .Q (new_AGEMA_signal_20908) ) ;
    buf_clk new_AGEMA_reg_buffer_8187 ( .C (clk), .D (new_AGEMA_signal_20910), .Q (new_AGEMA_signal_20911) ) ;
    buf_clk new_AGEMA_reg_buffer_8190 ( .C (clk), .D (new_AGEMA_signal_20913), .Q (new_AGEMA_signal_20914) ) ;
    buf_clk new_AGEMA_reg_buffer_8193 ( .C (clk), .D (new_AGEMA_signal_20916), .Q (new_AGEMA_signal_20917) ) ;
    buf_clk new_AGEMA_reg_buffer_8196 ( .C (clk), .D (new_AGEMA_signal_20919), .Q (new_AGEMA_signal_20920) ) ;
    buf_clk new_AGEMA_reg_buffer_8199 ( .C (clk), .D (new_AGEMA_signal_20922), .Q (new_AGEMA_signal_20923) ) ;
    buf_clk new_AGEMA_reg_buffer_8202 ( .C (clk), .D (new_AGEMA_signal_20925), .Q (new_AGEMA_signal_20926) ) ;
    buf_clk new_AGEMA_reg_buffer_8205 ( .C (clk), .D (new_AGEMA_signal_20928), .Q (new_AGEMA_signal_20929) ) ;
    buf_clk new_AGEMA_reg_buffer_8208 ( .C (clk), .D (new_AGEMA_signal_20931), .Q (new_AGEMA_signal_20932) ) ;
    buf_clk new_AGEMA_reg_buffer_8211 ( .C (clk), .D (new_AGEMA_signal_20934), .Q (new_AGEMA_signal_20935) ) ;
    buf_clk new_AGEMA_reg_buffer_8214 ( .C (clk), .D (new_AGEMA_signal_20937), .Q (new_AGEMA_signal_20938) ) ;
    buf_clk new_AGEMA_reg_buffer_8217 ( .C (clk), .D (new_AGEMA_signal_20940), .Q (new_AGEMA_signal_20941) ) ;
    buf_clk new_AGEMA_reg_buffer_8220 ( .C (clk), .D (new_AGEMA_signal_20943), .Q (new_AGEMA_signal_20944) ) ;
    buf_clk new_AGEMA_reg_buffer_8223 ( .C (clk), .D (new_AGEMA_signal_20946), .Q (new_AGEMA_signal_20947) ) ;
    buf_clk new_AGEMA_reg_buffer_8226 ( .C (clk), .D (new_AGEMA_signal_20949), .Q (new_AGEMA_signal_20950) ) ;
    buf_clk new_AGEMA_reg_buffer_8229 ( .C (clk), .D (new_AGEMA_signal_20952), .Q (new_AGEMA_signal_20953) ) ;
    buf_clk new_AGEMA_reg_buffer_8232 ( .C (clk), .D (new_AGEMA_signal_20955), .Q (new_AGEMA_signal_20956) ) ;
    buf_clk new_AGEMA_reg_buffer_8235 ( .C (clk), .D (new_AGEMA_signal_20958), .Q (new_AGEMA_signal_20959) ) ;
    buf_clk new_AGEMA_reg_buffer_8238 ( .C (clk), .D (new_AGEMA_signal_20961), .Q (new_AGEMA_signal_20962) ) ;
    buf_clk new_AGEMA_reg_buffer_8241 ( .C (clk), .D (new_AGEMA_signal_20964), .Q (new_AGEMA_signal_20965) ) ;
    buf_clk new_AGEMA_reg_buffer_8244 ( .C (clk), .D (new_AGEMA_signal_20967), .Q (new_AGEMA_signal_20968) ) ;
    buf_clk new_AGEMA_reg_buffer_8247 ( .C (clk), .D (new_AGEMA_signal_20970), .Q (new_AGEMA_signal_20971) ) ;
    buf_clk new_AGEMA_reg_buffer_8250 ( .C (clk), .D (new_AGEMA_signal_20973), .Q (new_AGEMA_signal_20974) ) ;
    buf_clk new_AGEMA_reg_buffer_8253 ( .C (clk), .D (new_AGEMA_signal_20976), .Q (new_AGEMA_signal_20977) ) ;
    buf_clk new_AGEMA_reg_buffer_8256 ( .C (clk), .D (new_AGEMA_signal_20979), .Q (new_AGEMA_signal_20980) ) ;
    buf_clk new_AGEMA_reg_buffer_8259 ( .C (clk), .D (new_AGEMA_signal_20982), .Q (new_AGEMA_signal_20983) ) ;
    buf_clk new_AGEMA_reg_buffer_8262 ( .C (clk), .D (new_AGEMA_signal_20985), .Q (new_AGEMA_signal_20986) ) ;
    buf_clk new_AGEMA_reg_buffer_8265 ( .C (clk), .D (new_AGEMA_signal_20988), .Q (new_AGEMA_signal_20989) ) ;
    buf_clk new_AGEMA_reg_buffer_8268 ( .C (clk), .D (new_AGEMA_signal_20991), .Q (new_AGEMA_signal_20992) ) ;
    buf_clk new_AGEMA_reg_buffer_8271 ( .C (clk), .D (new_AGEMA_signal_20994), .Q (new_AGEMA_signal_20995) ) ;
    buf_clk new_AGEMA_reg_buffer_8274 ( .C (clk), .D (new_AGEMA_signal_20997), .Q (new_AGEMA_signal_20998) ) ;
    buf_clk new_AGEMA_reg_buffer_8277 ( .C (clk), .D (new_AGEMA_signal_21000), .Q (new_AGEMA_signal_21001) ) ;
    buf_clk new_AGEMA_reg_buffer_8280 ( .C (clk), .D (new_AGEMA_signal_21003), .Q (new_AGEMA_signal_21004) ) ;
    buf_clk new_AGEMA_reg_buffer_8283 ( .C (clk), .D (new_AGEMA_signal_21006), .Q (new_AGEMA_signal_21007) ) ;
    buf_clk new_AGEMA_reg_buffer_8286 ( .C (clk), .D (new_AGEMA_signal_21009), .Q (new_AGEMA_signal_21010) ) ;
    buf_clk new_AGEMA_reg_buffer_8289 ( .C (clk), .D (new_AGEMA_signal_21012), .Q (new_AGEMA_signal_21013) ) ;
    buf_clk new_AGEMA_reg_buffer_8292 ( .C (clk), .D (new_AGEMA_signal_21015), .Q (new_AGEMA_signal_21016) ) ;
    buf_clk new_AGEMA_reg_buffer_8295 ( .C (clk), .D (new_AGEMA_signal_21018), .Q (new_AGEMA_signal_21019) ) ;
    buf_clk new_AGEMA_reg_buffer_8298 ( .C (clk), .D (new_AGEMA_signal_21021), .Q (new_AGEMA_signal_21022) ) ;
    buf_clk new_AGEMA_reg_buffer_8301 ( .C (clk), .D (new_AGEMA_signal_21024), .Q (new_AGEMA_signal_21025) ) ;
    buf_clk new_AGEMA_reg_buffer_8304 ( .C (clk), .D (new_AGEMA_signal_21027), .Q (new_AGEMA_signal_21028) ) ;
    buf_clk new_AGEMA_reg_buffer_8307 ( .C (clk), .D (new_AGEMA_signal_21030), .Q (new_AGEMA_signal_21031) ) ;
    buf_clk new_AGEMA_reg_buffer_8310 ( .C (clk), .D (new_AGEMA_signal_21033), .Q (new_AGEMA_signal_21034) ) ;
    buf_clk new_AGEMA_reg_buffer_8313 ( .C (clk), .D (new_AGEMA_signal_21036), .Q (new_AGEMA_signal_21037) ) ;
    buf_clk new_AGEMA_reg_buffer_8316 ( .C (clk), .D (new_AGEMA_signal_21039), .Q (new_AGEMA_signal_21040) ) ;
    buf_clk new_AGEMA_reg_buffer_8319 ( .C (clk), .D (new_AGEMA_signal_21042), .Q (new_AGEMA_signal_21043) ) ;
    buf_clk new_AGEMA_reg_buffer_8322 ( .C (clk), .D (new_AGEMA_signal_21045), .Q (new_AGEMA_signal_21046) ) ;
    buf_clk new_AGEMA_reg_buffer_8325 ( .C (clk), .D (new_AGEMA_signal_21048), .Q (new_AGEMA_signal_21049) ) ;
    buf_clk new_AGEMA_reg_buffer_8328 ( .C (clk), .D (new_AGEMA_signal_21051), .Q (new_AGEMA_signal_21052) ) ;
    buf_clk new_AGEMA_reg_buffer_8331 ( .C (clk), .D (new_AGEMA_signal_21054), .Q (new_AGEMA_signal_21055) ) ;
    buf_clk new_AGEMA_reg_buffer_8334 ( .C (clk), .D (new_AGEMA_signal_21057), .Q (new_AGEMA_signal_21058) ) ;
    buf_clk new_AGEMA_reg_buffer_8337 ( .C (clk), .D (new_AGEMA_signal_21060), .Q (new_AGEMA_signal_21061) ) ;
    buf_clk new_AGEMA_reg_buffer_8340 ( .C (clk), .D (new_AGEMA_signal_21063), .Q (new_AGEMA_signal_21064) ) ;
    buf_clk new_AGEMA_reg_buffer_8343 ( .C (clk), .D (new_AGEMA_signal_21066), .Q (new_AGEMA_signal_21067) ) ;
    buf_clk new_AGEMA_reg_buffer_8346 ( .C (clk), .D (new_AGEMA_signal_21069), .Q (new_AGEMA_signal_21070) ) ;
    buf_clk new_AGEMA_reg_buffer_8349 ( .C (clk), .D (new_AGEMA_signal_21072), .Q (new_AGEMA_signal_21073) ) ;
    buf_clk new_AGEMA_reg_buffer_8352 ( .C (clk), .D (new_AGEMA_signal_21075), .Q (new_AGEMA_signal_21076) ) ;
    buf_clk new_AGEMA_reg_buffer_8355 ( .C (clk), .D (new_AGEMA_signal_21078), .Q (new_AGEMA_signal_21079) ) ;
    buf_clk new_AGEMA_reg_buffer_8358 ( .C (clk), .D (new_AGEMA_signal_21081), .Q (new_AGEMA_signal_21082) ) ;
    buf_clk new_AGEMA_reg_buffer_8361 ( .C (clk), .D (new_AGEMA_signal_21084), .Q (new_AGEMA_signal_21085) ) ;
    buf_clk new_AGEMA_reg_buffer_8364 ( .C (clk), .D (new_AGEMA_signal_21087), .Q (new_AGEMA_signal_21088) ) ;
    buf_clk new_AGEMA_reg_buffer_8367 ( .C (clk), .D (new_AGEMA_signal_21090), .Q (new_AGEMA_signal_21091) ) ;
    buf_clk new_AGEMA_reg_buffer_8370 ( .C (clk), .D (new_AGEMA_signal_21093), .Q (new_AGEMA_signal_21094) ) ;
    buf_clk new_AGEMA_reg_buffer_8373 ( .C (clk), .D (new_AGEMA_signal_21096), .Q (new_AGEMA_signal_21097) ) ;
    buf_clk new_AGEMA_reg_buffer_8376 ( .C (clk), .D (new_AGEMA_signal_21099), .Q (new_AGEMA_signal_21100) ) ;
    buf_clk new_AGEMA_reg_buffer_8379 ( .C (clk), .D (new_AGEMA_signal_21102), .Q (new_AGEMA_signal_21103) ) ;
    buf_clk new_AGEMA_reg_buffer_8382 ( .C (clk), .D (new_AGEMA_signal_21105), .Q (new_AGEMA_signal_21106) ) ;
    buf_clk new_AGEMA_reg_buffer_8385 ( .C (clk), .D (new_AGEMA_signal_21108), .Q (new_AGEMA_signal_21109) ) ;
    buf_clk new_AGEMA_reg_buffer_8388 ( .C (clk), .D (new_AGEMA_signal_21111), .Q (new_AGEMA_signal_21112) ) ;
    buf_clk new_AGEMA_reg_buffer_8391 ( .C (clk), .D (new_AGEMA_signal_21114), .Q (new_AGEMA_signal_21115) ) ;
    buf_clk new_AGEMA_reg_buffer_8394 ( .C (clk), .D (new_AGEMA_signal_21117), .Q (new_AGEMA_signal_21118) ) ;
    buf_clk new_AGEMA_reg_buffer_8397 ( .C (clk), .D (new_AGEMA_signal_21120), .Q (new_AGEMA_signal_21121) ) ;
    buf_clk new_AGEMA_reg_buffer_8400 ( .C (clk), .D (new_AGEMA_signal_21123), .Q (new_AGEMA_signal_21124) ) ;
    buf_clk new_AGEMA_reg_buffer_8403 ( .C (clk), .D (new_AGEMA_signal_21126), .Q (new_AGEMA_signal_21127) ) ;
    buf_clk new_AGEMA_reg_buffer_8406 ( .C (clk), .D (new_AGEMA_signal_21129), .Q (new_AGEMA_signal_21130) ) ;
    buf_clk new_AGEMA_reg_buffer_8409 ( .C (clk), .D (new_AGEMA_signal_21132), .Q (new_AGEMA_signal_21133) ) ;
    buf_clk new_AGEMA_reg_buffer_8412 ( .C (clk), .D (new_AGEMA_signal_21135), .Q (new_AGEMA_signal_21136) ) ;
    buf_clk new_AGEMA_reg_buffer_8415 ( .C (clk), .D (new_AGEMA_signal_21138), .Q (new_AGEMA_signal_21139) ) ;
    buf_clk new_AGEMA_reg_buffer_8418 ( .C (clk), .D (new_AGEMA_signal_21141), .Q (new_AGEMA_signal_21142) ) ;
    buf_clk new_AGEMA_reg_buffer_8421 ( .C (clk), .D (new_AGEMA_signal_21144), .Q (new_AGEMA_signal_21145) ) ;
    buf_clk new_AGEMA_reg_buffer_8424 ( .C (clk), .D (new_AGEMA_signal_21147), .Q (new_AGEMA_signal_21148) ) ;
    buf_clk new_AGEMA_reg_buffer_8427 ( .C (clk), .D (new_AGEMA_signal_21150), .Q (new_AGEMA_signal_21151) ) ;
    buf_clk new_AGEMA_reg_buffer_8430 ( .C (clk), .D (new_AGEMA_signal_21153), .Q (new_AGEMA_signal_21154) ) ;
    buf_clk new_AGEMA_reg_buffer_8433 ( .C (clk), .D (new_AGEMA_signal_21156), .Q (new_AGEMA_signal_21157) ) ;
    buf_clk new_AGEMA_reg_buffer_8436 ( .C (clk), .D (new_AGEMA_signal_21159), .Q (new_AGEMA_signal_21160) ) ;
    buf_clk new_AGEMA_reg_buffer_8439 ( .C (clk), .D (new_AGEMA_signal_21162), .Q (new_AGEMA_signal_21163) ) ;
    buf_clk new_AGEMA_reg_buffer_8442 ( .C (clk), .D (new_AGEMA_signal_21165), .Q (new_AGEMA_signal_21166) ) ;
    buf_clk new_AGEMA_reg_buffer_8445 ( .C (clk), .D (new_AGEMA_signal_21168), .Q (new_AGEMA_signal_21169) ) ;
    buf_clk new_AGEMA_reg_buffer_8448 ( .C (clk), .D (new_AGEMA_signal_21171), .Q (new_AGEMA_signal_21172) ) ;
    buf_clk new_AGEMA_reg_buffer_8451 ( .C (clk), .D (new_AGEMA_signal_21174), .Q (new_AGEMA_signal_21175) ) ;
    buf_clk new_AGEMA_reg_buffer_8454 ( .C (clk), .D (new_AGEMA_signal_21177), .Q (new_AGEMA_signal_21178) ) ;
    buf_clk new_AGEMA_reg_buffer_8457 ( .C (clk), .D (new_AGEMA_signal_21180), .Q (new_AGEMA_signal_21181) ) ;
    buf_clk new_AGEMA_reg_buffer_8460 ( .C (clk), .D (new_AGEMA_signal_21183), .Q (new_AGEMA_signal_21184) ) ;
    buf_clk new_AGEMA_reg_buffer_8463 ( .C (clk), .D (new_AGEMA_signal_21186), .Q (new_AGEMA_signal_21187) ) ;
    buf_clk new_AGEMA_reg_buffer_8466 ( .C (clk), .D (new_AGEMA_signal_21189), .Q (new_AGEMA_signal_21190) ) ;
    buf_clk new_AGEMA_reg_buffer_8469 ( .C (clk), .D (new_AGEMA_signal_21192), .Q (new_AGEMA_signal_21193) ) ;
    buf_clk new_AGEMA_reg_buffer_8472 ( .C (clk), .D (new_AGEMA_signal_21195), .Q (new_AGEMA_signal_21196) ) ;
    buf_clk new_AGEMA_reg_buffer_8475 ( .C (clk), .D (new_AGEMA_signal_21198), .Q (new_AGEMA_signal_21199) ) ;
    buf_clk new_AGEMA_reg_buffer_8478 ( .C (clk), .D (new_AGEMA_signal_21201), .Q (new_AGEMA_signal_21202) ) ;
    buf_clk new_AGEMA_reg_buffer_8481 ( .C (clk), .D (new_AGEMA_signal_21204), .Q (new_AGEMA_signal_21205) ) ;
    buf_clk new_AGEMA_reg_buffer_8484 ( .C (clk), .D (new_AGEMA_signal_21207), .Q (new_AGEMA_signal_21208) ) ;
    buf_clk new_AGEMA_reg_buffer_8487 ( .C (clk), .D (new_AGEMA_signal_21210), .Q (new_AGEMA_signal_21211) ) ;
    buf_clk new_AGEMA_reg_buffer_8490 ( .C (clk), .D (new_AGEMA_signal_21213), .Q (new_AGEMA_signal_21214) ) ;
    buf_clk new_AGEMA_reg_buffer_8493 ( .C (clk), .D (new_AGEMA_signal_21216), .Q (new_AGEMA_signal_21217) ) ;
    buf_clk new_AGEMA_reg_buffer_8496 ( .C (clk), .D (new_AGEMA_signal_21219), .Q (new_AGEMA_signal_21220) ) ;
    buf_clk new_AGEMA_reg_buffer_8499 ( .C (clk), .D (new_AGEMA_signal_21222), .Q (new_AGEMA_signal_21223) ) ;
    buf_clk new_AGEMA_reg_buffer_8502 ( .C (clk), .D (new_AGEMA_signal_21225), .Q (new_AGEMA_signal_21226) ) ;
    buf_clk new_AGEMA_reg_buffer_8505 ( .C (clk), .D (new_AGEMA_signal_21228), .Q (new_AGEMA_signal_21229) ) ;
    buf_clk new_AGEMA_reg_buffer_8508 ( .C (clk), .D (new_AGEMA_signal_21231), .Q (new_AGEMA_signal_21232) ) ;
    buf_clk new_AGEMA_reg_buffer_8511 ( .C (clk), .D (new_AGEMA_signal_21234), .Q (new_AGEMA_signal_21235) ) ;
    buf_clk new_AGEMA_reg_buffer_8514 ( .C (clk), .D (new_AGEMA_signal_21237), .Q (new_AGEMA_signal_21238) ) ;
    buf_clk new_AGEMA_reg_buffer_8517 ( .C (clk), .D (new_AGEMA_signal_21240), .Q (new_AGEMA_signal_21241) ) ;
    buf_clk new_AGEMA_reg_buffer_8520 ( .C (clk), .D (new_AGEMA_signal_21243), .Q (new_AGEMA_signal_21244) ) ;
    buf_clk new_AGEMA_reg_buffer_8523 ( .C (clk), .D (new_AGEMA_signal_21246), .Q (new_AGEMA_signal_21247) ) ;
    buf_clk new_AGEMA_reg_buffer_8526 ( .C (clk), .D (new_AGEMA_signal_21249), .Q (new_AGEMA_signal_21250) ) ;
    buf_clk new_AGEMA_reg_buffer_8529 ( .C (clk), .D (new_AGEMA_signal_21252), .Q (new_AGEMA_signal_21253) ) ;
    buf_clk new_AGEMA_reg_buffer_8532 ( .C (clk), .D (new_AGEMA_signal_21255), .Q (new_AGEMA_signal_21256) ) ;
    buf_clk new_AGEMA_reg_buffer_8535 ( .C (clk), .D (new_AGEMA_signal_21258), .Q (new_AGEMA_signal_21259) ) ;
    buf_clk new_AGEMA_reg_buffer_8538 ( .C (clk), .D (new_AGEMA_signal_21261), .Q (new_AGEMA_signal_21262) ) ;
    buf_clk new_AGEMA_reg_buffer_8541 ( .C (clk), .D (new_AGEMA_signal_21264), .Q (new_AGEMA_signal_21265) ) ;
    buf_clk new_AGEMA_reg_buffer_8544 ( .C (clk), .D (new_AGEMA_signal_21267), .Q (new_AGEMA_signal_21268) ) ;
    buf_clk new_AGEMA_reg_buffer_8547 ( .C (clk), .D (new_AGEMA_signal_21270), .Q (new_AGEMA_signal_21271) ) ;
    buf_clk new_AGEMA_reg_buffer_8550 ( .C (clk), .D (new_AGEMA_signal_21273), .Q (new_AGEMA_signal_21274) ) ;
    buf_clk new_AGEMA_reg_buffer_8553 ( .C (clk), .D (new_AGEMA_signal_21276), .Q (new_AGEMA_signal_21277) ) ;
    buf_clk new_AGEMA_reg_buffer_8556 ( .C (clk), .D (new_AGEMA_signal_21279), .Q (new_AGEMA_signal_21280) ) ;
    buf_clk new_AGEMA_reg_buffer_8559 ( .C (clk), .D (new_AGEMA_signal_21282), .Q (new_AGEMA_signal_21283) ) ;
    buf_clk new_AGEMA_reg_buffer_8562 ( .C (clk), .D (new_AGEMA_signal_21285), .Q (new_AGEMA_signal_21286) ) ;
    buf_clk new_AGEMA_reg_buffer_8565 ( .C (clk), .D (new_AGEMA_signal_21288), .Q (new_AGEMA_signal_21289) ) ;
    buf_clk new_AGEMA_reg_buffer_8568 ( .C (clk), .D (new_AGEMA_signal_21291), .Q (new_AGEMA_signal_21292) ) ;
    buf_clk new_AGEMA_reg_buffer_8571 ( .C (clk), .D (new_AGEMA_signal_21294), .Q (new_AGEMA_signal_21295) ) ;
    buf_clk new_AGEMA_reg_buffer_8574 ( .C (clk), .D (new_AGEMA_signal_21297), .Q (new_AGEMA_signal_21298) ) ;
    buf_clk new_AGEMA_reg_buffer_8577 ( .C (clk), .D (new_AGEMA_signal_21300), .Q (new_AGEMA_signal_21301) ) ;
    buf_clk new_AGEMA_reg_buffer_8580 ( .C (clk), .D (new_AGEMA_signal_21303), .Q (new_AGEMA_signal_21304) ) ;
    buf_clk new_AGEMA_reg_buffer_8583 ( .C (clk), .D (new_AGEMA_signal_21306), .Q (new_AGEMA_signal_21307) ) ;
    buf_clk new_AGEMA_reg_buffer_8586 ( .C (clk), .D (new_AGEMA_signal_21309), .Q (new_AGEMA_signal_21310) ) ;
    buf_clk new_AGEMA_reg_buffer_8589 ( .C (clk), .D (new_AGEMA_signal_21312), .Q (new_AGEMA_signal_21313) ) ;
    buf_clk new_AGEMA_reg_buffer_8592 ( .C (clk), .D (new_AGEMA_signal_21315), .Q (new_AGEMA_signal_21316) ) ;
    buf_clk new_AGEMA_reg_buffer_8595 ( .C (clk), .D (new_AGEMA_signal_21318), .Q (new_AGEMA_signal_21319) ) ;
    buf_clk new_AGEMA_reg_buffer_8598 ( .C (clk), .D (new_AGEMA_signal_21321), .Q (new_AGEMA_signal_21322) ) ;
    buf_clk new_AGEMA_reg_buffer_8601 ( .C (clk), .D (new_AGEMA_signal_21324), .Q (new_AGEMA_signal_21325) ) ;
    buf_clk new_AGEMA_reg_buffer_8604 ( .C (clk), .D (new_AGEMA_signal_21327), .Q (new_AGEMA_signal_21328) ) ;
    buf_clk new_AGEMA_reg_buffer_8607 ( .C (clk), .D (new_AGEMA_signal_21330), .Q (new_AGEMA_signal_21331) ) ;
    buf_clk new_AGEMA_reg_buffer_8610 ( .C (clk), .D (new_AGEMA_signal_21333), .Q (new_AGEMA_signal_21334) ) ;
    buf_clk new_AGEMA_reg_buffer_8613 ( .C (clk), .D (new_AGEMA_signal_21336), .Q (new_AGEMA_signal_21337) ) ;
    buf_clk new_AGEMA_reg_buffer_8616 ( .C (clk), .D (new_AGEMA_signal_21339), .Q (new_AGEMA_signal_21340) ) ;
    buf_clk new_AGEMA_reg_buffer_8619 ( .C (clk), .D (new_AGEMA_signal_21342), .Q (new_AGEMA_signal_21343) ) ;
    buf_clk new_AGEMA_reg_buffer_8622 ( .C (clk), .D (new_AGEMA_signal_21345), .Q (new_AGEMA_signal_21346) ) ;
    buf_clk new_AGEMA_reg_buffer_8625 ( .C (clk), .D (new_AGEMA_signal_21348), .Q (new_AGEMA_signal_21349) ) ;
    buf_clk new_AGEMA_reg_buffer_8628 ( .C (clk), .D (new_AGEMA_signal_21351), .Q (new_AGEMA_signal_21352) ) ;
    buf_clk new_AGEMA_reg_buffer_8631 ( .C (clk), .D (new_AGEMA_signal_21354), .Q (new_AGEMA_signal_21355) ) ;
    buf_clk new_AGEMA_reg_buffer_8634 ( .C (clk), .D (new_AGEMA_signal_21357), .Q (new_AGEMA_signal_21358) ) ;
    buf_clk new_AGEMA_reg_buffer_8637 ( .C (clk), .D (new_AGEMA_signal_21360), .Q (new_AGEMA_signal_21361) ) ;
    buf_clk new_AGEMA_reg_buffer_8640 ( .C (clk), .D (new_AGEMA_signal_21363), .Q (new_AGEMA_signal_21364) ) ;
    buf_clk new_AGEMA_reg_buffer_8643 ( .C (clk), .D (new_AGEMA_signal_21366), .Q (new_AGEMA_signal_21367) ) ;
    buf_clk new_AGEMA_reg_buffer_8646 ( .C (clk), .D (new_AGEMA_signal_21369), .Q (new_AGEMA_signal_21370) ) ;
    buf_clk new_AGEMA_reg_buffer_8649 ( .C (clk), .D (new_AGEMA_signal_21372), .Q (new_AGEMA_signal_21373) ) ;
    buf_clk new_AGEMA_reg_buffer_8652 ( .C (clk), .D (new_AGEMA_signal_21375), .Q (new_AGEMA_signal_21376) ) ;
    buf_clk new_AGEMA_reg_buffer_8655 ( .C (clk), .D (new_AGEMA_signal_21378), .Q (new_AGEMA_signal_21379) ) ;
    buf_clk new_AGEMA_reg_buffer_8658 ( .C (clk), .D (new_AGEMA_signal_21381), .Q (new_AGEMA_signal_21382) ) ;
    buf_clk new_AGEMA_reg_buffer_8661 ( .C (clk), .D (new_AGEMA_signal_21384), .Q (new_AGEMA_signal_21385) ) ;
    buf_clk new_AGEMA_reg_buffer_8664 ( .C (clk), .D (new_AGEMA_signal_21387), .Q (new_AGEMA_signal_21388) ) ;
    buf_clk new_AGEMA_reg_buffer_8667 ( .C (clk), .D (new_AGEMA_signal_21390), .Q (new_AGEMA_signal_21391) ) ;
    buf_clk new_AGEMA_reg_buffer_8670 ( .C (clk), .D (new_AGEMA_signal_21393), .Q (new_AGEMA_signal_21394) ) ;
    buf_clk new_AGEMA_reg_buffer_8673 ( .C (clk), .D (new_AGEMA_signal_21396), .Q (new_AGEMA_signal_21397) ) ;
    buf_clk new_AGEMA_reg_buffer_8676 ( .C (clk), .D (new_AGEMA_signal_21399), .Q (new_AGEMA_signal_21400) ) ;
    buf_clk new_AGEMA_reg_buffer_8679 ( .C (clk), .D (new_AGEMA_signal_21402), .Q (new_AGEMA_signal_21403) ) ;
    buf_clk new_AGEMA_reg_buffer_8682 ( .C (clk), .D (new_AGEMA_signal_21405), .Q (new_AGEMA_signal_21406) ) ;
    buf_clk new_AGEMA_reg_buffer_8685 ( .C (clk), .D (new_AGEMA_signal_21408), .Q (new_AGEMA_signal_21409) ) ;
    buf_clk new_AGEMA_reg_buffer_8688 ( .C (clk), .D (new_AGEMA_signal_21411), .Q (new_AGEMA_signal_21412) ) ;
    buf_clk new_AGEMA_reg_buffer_8691 ( .C (clk), .D (new_AGEMA_signal_21414), .Q (new_AGEMA_signal_21415) ) ;
    buf_clk new_AGEMA_reg_buffer_8694 ( .C (clk), .D (new_AGEMA_signal_21417), .Q (new_AGEMA_signal_21418) ) ;
    buf_clk new_AGEMA_reg_buffer_8697 ( .C (clk), .D (new_AGEMA_signal_21420), .Q (new_AGEMA_signal_21421) ) ;
    buf_clk new_AGEMA_reg_buffer_8700 ( .C (clk), .D (new_AGEMA_signal_21423), .Q (new_AGEMA_signal_21424) ) ;
    buf_clk new_AGEMA_reg_buffer_8703 ( .C (clk), .D (new_AGEMA_signal_21426), .Q (new_AGEMA_signal_21427) ) ;
    buf_clk new_AGEMA_reg_buffer_8706 ( .C (clk), .D (new_AGEMA_signal_21429), .Q (new_AGEMA_signal_21430) ) ;
    buf_clk new_AGEMA_reg_buffer_8709 ( .C (clk), .D (new_AGEMA_signal_21432), .Q (new_AGEMA_signal_21433) ) ;
    buf_clk new_AGEMA_reg_buffer_8712 ( .C (clk), .D (new_AGEMA_signal_21435), .Q (new_AGEMA_signal_21436) ) ;
    buf_clk new_AGEMA_reg_buffer_8715 ( .C (clk), .D (new_AGEMA_signal_21438), .Q (new_AGEMA_signal_21439) ) ;
    buf_clk new_AGEMA_reg_buffer_8718 ( .C (clk), .D (new_AGEMA_signal_21441), .Q (new_AGEMA_signal_21442) ) ;
    buf_clk new_AGEMA_reg_buffer_8721 ( .C (clk), .D (new_AGEMA_signal_21444), .Q (new_AGEMA_signal_21445) ) ;
    buf_clk new_AGEMA_reg_buffer_8724 ( .C (clk), .D (new_AGEMA_signal_21447), .Q (new_AGEMA_signal_21448) ) ;
    buf_clk new_AGEMA_reg_buffer_8727 ( .C (clk), .D (new_AGEMA_signal_21450), .Q (new_AGEMA_signal_21451) ) ;
    buf_clk new_AGEMA_reg_buffer_8730 ( .C (clk), .D (new_AGEMA_signal_21453), .Q (new_AGEMA_signal_21454) ) ;
    buf_clk new_AGEMA_reg_buffer_8733 ( .C (clk), .D (new_AGEMA_signal_21456), .Q (new_AGEMA_signal_21457) ) ;
    buf_clk new_AGEMA_reg_buffer_8736 ( .C (clk), .D (new_AGEMA_signal_21459), .Q (new_AGEMA_signal_21460) ) ;
    buf_clk new_AGEMA_reg_buffer_8739 ( .C (clk), .D (new_AGEMA_signal_21462), .Q (new_AGEMA_signal_21463) ) ;
    buf_clk new_AGEMA_reg_buffer_8742 ( .C (clk), .D (new_AGEMA_signal_21465), .Q (new_AGEMA_signal_21466) ) ;
    buf_clk new_AGEMA_reg_buffer_8745 ( .C (clk), .D (new_AGEMA_signal_21468), .Q (new_AGEMA_signal_21469) ) ;
    buf_clk new_AGEMA_reg_buffer_8748 ( .C (clk), .D (new_AGEMA_signal_21471), .Q (new_AGEMA_signal_21472) ) ;
    buf_clk new_AGEMA_reg_buffer_8751 ( .C (clk), .D (new_AGEMA_signal_21474), .Q (new_AGEMA_signal_21475) ) ;
    buf_clk new_AGEMA_reg_buffer_8754 ( .C (clk), .D (new_AGEMA_signal_21477), .Q (new_AGEMA_signal_21478) ) ;
    buf_clk new_AGEMA_reg_buffer_8757 ( .C (clk), .D (new_AGEMA_signal_21480), .Q (new_AGEMA_signal_21481) ) ;
    buf_clk new_AGEMA_reg_buffer_8760 ( .C (clk), .D (new_AGEMA_signal_21483), .Q (new_AGEMA_signal_21484) ) ;
    buf_clk new_AGEMA_reg_buffer_8763 ( .C (clk), .D (new_AGEMA_signal_21486), .Q (new_AGEMA_signal_21487) ) ;
    buf_clk new_AGEMA_reg_buffer_8766 ( .C (clk), .D (new_AGEMA_signal_21489), .Q (new_AGEMA_signal_21490) ) ;
    buf_clk new_AGEMA_reg_buffer_8769 ( .C (clk), .D (new_AGEMA_signal_21492), .Q (new_AGEMA_signal_21493) ) ;
    buf_clk new_AGEMA_reg_buffer_8772 ( .C (clk), .D (new_AGEMA_signal_21495), .Q (new_AGEMA_signal_21496) ) ;
    buf_clk new_AGEMA_reg_buffer_8775 ( .C (clk), .D (new_AGEMA_signal_21498), .Q (new_AGEMA_signal_21499) ) ;
    buf_clk new_AGEMA_reg_buffer_8778 ( .C (clk), .D (new_AGEMA_signal_21501), .Q (new_AGEMA_signal_21502) ) ;
    buf_clk new_AGEMA_reg_buffer_8781 ( .C (clk), .D (new_AGEMA_signal_21504), .Q (new_AGEMA_signal_21505) ) ;
    buf_clk new_AGEMA_reg_buffer_8784 ( .C (clk), .D (new_AGEMA_signal_21507), .Q (new_AGEMA_signal_21508) ) ;
    buf_clk new_AGEMA_reg_buffer_8787 ( .C (clk), .D (new_AGEMA_signal_21510), .Q (new_AGEMA_signal_21511) ) ;
    buf_clk new_AGEMA_reg_buffer_8790 ( .C (clk), .D (new_AGEMA_signal_21513), .Q (new_AGEMA_signal_21514) ) ;
    buf_clk new_AGEMA_reg_buffer_8793 ( .C (clk), .D (new_AGEMA_signal_21516), .Q (new_AGEMA_signal_21517) ) ;
    buf_clk new_AGEMA_reg_buffer_8796 ( .C (clk), .D (new_AGEMA_signal_21519), .Q (new_AGEMA_signal_21520) ) ;
    buf_clk new_AGEMA_reg_buffer_8799 ( .C (clk), .D (new_AGEMA_signal_21522), .Q (new_AGEMA_signal_21523) ) ;
    buf_clk new_AGEMA_reg_buffer_8802 ( .C (clk), .D (new_AGEMA_signal_21525), .Q (new_AGEMA_signal_21526) ) ;
    buf_clk new_AGEMA_reg_buffer_8805 ( .C (clk), .D (new_AGEMA_signal_21528), .Q (new_AGEMA_signal_21529) ) ;
    buf_clk new_AGEMA_reg_buffer_8808 ( .C (clk), .D (new_AGEMA_signal_21531), .Q (new_AGEMA_signal_21532) ) ;
    buf_clk new_AGEMA_reg_buffer_8811 ( .C (clk), .D (new_AGEMA_signal_21534), .Q (new_AGEMA_signal_21535) ) ;
    buf_clk new_AGEMA_reg_buffer_8814 ( .C (clk), .D (new_AGEMA_signal_21537), .Q (new_AGEMA_signal_21538) ) ;
    buf_clk new_AGEMA_reg_buffer_8817 ( .C (clk), .D (new_AGEMA_signal_21540), .Q (new_AGEMA_signal_21541) ) ;
    buf_clk new_AGEMA_reg_buffer_8820 ( .C (clk), .D (new_AGEMA_signal_21543), .Q (new_AGEMA_signal_21544) ) ;
    buf_clk new_AGEMA_reg_buffer_8823 ( .C (clk), .D (new_AGEMA_signal_21546), .Q (new_AGEMA_signal_21547) ) ;
    buf_clk new_AGEMA_reg_buffer_8826 ( .C (clk), .D (new_AGEMA_signal_21549), .Q (new_AGEMA_signal_21550) ) ;
    buf_clk new_AGEMA_reg_buffer_8829 ( .C (clk), .D (new_AGEMA_signal_21552), .Q (new_AGEMA_signal_21553) ) ;
    buf_clk new_AGEMA_reg_buffer_8832 ( .C (clk), .D (new_AGEMA_signal_21555), .Q (new_AGEMA_signal_21556) ) ;
    buf_clk new_AGEMA_reg_buffer_8835 ( .C (clk), .D (new_AGEMA_signal_21558), .Q (new_AGEMA_signal_21559) ) ;
    buf_clk new_AGEMA_reg_buffer_8838 ( .C (clk), .D (new_AGEMA_signal_21561), .Q (new_AGEMA_signal_21562) ) ;
    buf_clk new_AGEMA_reg_buffer_8841 ( .C (clk), .D (new_AGEMA_signal_21564), .Q (new_AGEMA_signal_21565) ) ;
    buf_clk new_AGEMA_reg_buffer_8844 ( .C (clk), .D (new_AGEMA_signal_21567), .Q (new_AGEMA_signal_21568) ) ;
    buf_clk new_AGEMA_reg_buffer_8847 ( .C (clk), .D (new_AGEMA_signal_21570), .Q (new_AGEMA_signal_21571) ) ;
    buf_clk new_AGEMA_reg_buffer_8850 ( .C (clk), .D (new_AGEMA_signal_21573), .Q (new_AGEMA_signal_21574) ) ;
    buf_clk new_AGEMA_reg_buffer_8853 ( .C (clk), .D (new_AGEMA_signal_21576), .Q (new_AGEMA_signal_21577) ) ;
    buf_clk new_AGEMA_reg_buffer_8856 ( .C (clk), .D (new_AGEMA_signal_21579), .Q (new_AGEMA_signal_21580) ) ;
    buf_clk new_AGEMA_reg_buffer_8859 ( .C (clk), .D (new_AGEMA_signal_21582), .Q (new_AGEMA_signal_21583) ) ;
    buf_clk new_AGEMA_reg_buffer_8862 ( .C (clk), .D (new_AGEMA_signal_21585), .Q (new_AGEMA_signal_21586) ) ;
    buf_clk new_AGEMA_reg_buffer_8865 ( .C (clk), .D (new_AGEMA_signal_21588), .Q (new_AGEMA_signal_21589) ) ;
    buf_clk new_AGEMA_reg_buffer_8868 ( .C (clk), .D (new_AGEMA_signal_21591), .Q (new_AGEMA_signal_21592) ) ;
    buf_clk new_AGEMA_reg_buffer_8871 ( .C (clk), .D (new_AGEMA_signal_21594), .Q (new_AGEMA_signal_21595) ) ;
    buf_clk new_AGEMA_reg_buffer_8874 ( .C (clk), .D (new_AGEMA_signal_21597), .Q (new_AGEMA_signal_21598) ) ;
    buf_clk new_AGEMA_reg_buffer_8877 ( .C (clk), .D (new_AGEMA_signal_21600), .Q (new_AGEMA_signal_21601) ) ;
    buf_clk new_AGEMA_reg_buffer_8880 ( .C (clk), .D (new_AGEMA_signal_21603), .Q (new_AGEMA_signal_21604) ) ;
    buf_clk new_AGEMA_reg_buffer_8883 ( .C (clk), .D (new_AGEMA_signal_21606), .Q (new_AGEMA_signal_21607) ) ;
    buf_clk new_AGEMA_reg_buffer_8886 ( .C (clk), .D (new_AGEMA_signal_21609), .Q (new_AGEMA_signal_21610) ) ;
    buf_clk new_AGEMA_reg_buffer_8889 ( .C (clk), .D (new_AGEMA_signal_21612), .Q (new_AGEMA_signal_21613) ) ;
    buf_clk new_AGEMA_reg_buffer_8892 ( .C (clk), .D (new_AGEMA_signal_21615), .Q (new_AGEMA_signal_21616) ) ;
    buf_clk new_AGEMA_reg_buffer_8895 ( .C (clk), .D (new_AGEMA_signal_21618), .Q (new_AGEMA_signal_21619) ) ;
    buf_clk new_AGEMA_reg_buffer_8898 ( .C (clk), .D (new_AGEMA_signal_21621), .Q (new_AGEMA_signal_21622) ) ;
    buf_clk new_AGEMA_reg_buffer_8901 ( .C (clk), .D (new_AGEMA_signal_21624), .Q (new_AGEMA_signal_21625) ) ;
    buf_clk new_AGEMA_reg_buffer_8904 ( .C (clk), .D (new_AGEMA_signal_21627), .Q (new_AGEMA_signal_21628) ) ;
    buf_clk new_AGEMA_reg_buffer_8907 ( .C (clk), .D (new_AGEMA_signal_21630), .Q (new_AGEMA_signal_21631) ) ;
    buf_clk new_AGEMA_reg_buffer_8910 ( .C (clk), .D (new_AGEMA_signal_21633), .Q (new_AGEMA_signal_21634) ) ;
    buf_clk new_AGEMA_reg_buffer_8913 ( .C (clk), .D (new_AGEMA_signal_21636), .Q (new_AGEMA_signal_21637) ) ;
    buf_clk new_AGEMA_reg_buffer_8916 ( .C (clk), .D (new_AGEMA_signal_21639), .Q (new_AGEMA_signal_21640) ) ;
    buf_clk new_AGEMA_reg_buffer_8919 ( .C (clk), .D (new_AGEMA_signal_21642), .Q (new_AGEMA_signal_21643) ) ;
    buf_clk new_AGEMA_reg_buffer_8922 ( .C (clk), .D (new_AGEMA_signal_21645), .Q (new_AGEMA_signal_21646) ) ;
    buf_clk new_AGEMA_reg_buffer_8925 ( .C (clk), .D (new_AGEMA_signal_21648), .Q (new_AGEMA_signal_21649) ) ;
    buf_clk new_AGEMA_reg_buffer_8928 ( .C (clk), .D (new_AGEMA_signal_21651), .Q (new_AGEMA_signal_21652) ) ;
    buf_clk new_AGEMA_reg_buffer_8931 ( .C (clk), .D (new_AGEMA_signal_21654), .Q (new_AGEMA_signal_21655) ) ;
    buf_clk new_AGEMA_reg_buffer_8934 ( .C (clk), .D (new_AGEMA_signal_21657), .Q (new_AGEMA_signal_21658) ) ;
    buf_clk new_AGEMA_reg_buffer_8937 ( .C (clk), .D (new_AGEMA_signal_21660), .Q (new_AGEMA_signal_21661) ) ;
    buf_clk new_AGEMA_reg_buffer_8940 ( .C (clk), .D (new_AGEMA_signal_21663), .Q (new_AGEMA_signal_21664) ) ;
    buf_clk new_AGEMA_reg_buffer_8943 ( .C (clk), .D (new_AGEMA_signal_21666), .Q (new_AGEMA_signal_21667) ) ;
    buf_clk new_AGEMA_reg_buffer_8946 ( .C (clk), .D (new_AGEMA_signal_21669), .Q (new_AGEMA_signal_21670) ) ;
    buf_clk new_AGEMA_reg_buffer_8949 ( .C (clk), .D (new_AGEMA_signal_21672), .Q (new_AGEMA_signal_21673) ) ;
    buf_clk new_AGEMA_reg_buffer_8952 ( .C (clk), .D (new_AGEMA_signal_21675), .Q (new_AGEMA_signal_21676) ) ;
    buf_clk new_AGEMA_reg_buffer_8955 ( .C (clk), .D (new_AGEMA_signal_21678), .Q (new_AGEMA_signal_21679) ) ;
    buf_clk new_AGEMA_reg_buffer_8958 ( .C (clk), .D (new_AGEMA_signal_21681), .Q (new_AGEMA_signal_21682) ) ;
    buf_clk new_AGEMA_reg_buffer_8961 ( .C (clk), .D (new_AGEMA_signal_21684), .Q (new_AGEMA_signal_21685) ) ;
    buf_clk new_AGEMA_reg_buffer_8964 ( .C (clk), .D (new_AGEMA_signal_21687), .Q (new_AGEMA_signal_21688) ) ;
    buf_clk new_AGEMA_reg_buffer_8967 ( .C (clk), .D (new_AGEMA_signal_21690), .Q (new_AGEMA_signal_21691) ) ;
    buf_clk new_AGEMA_reg_buffer_8970 ( .C (clk), .D (new_AGEMA_signal_21693), .Q (new_AGEMA_signal_21694) ) ;
    buf_clk new_AGEMA_reg_buffer_8973 ( .C (clk), .D (new_AGEMA_signal_21696), .Q (new_AGEMA_signal_21697) ) ;
    buf_clk new_AGEMA_reg_buffer_8976 ( .C (clk), .D (new_AGEMA_signal_21699), .Q (new_AGEMA_signal_21700) ) ;
    buf_clk new_AGEMA_reg_buffer_8979 ( .C (clk), .D (new_AGEMA_signal_21702), .Q (new_AGEMA_signal_21703) ) ;
    buf_clk new_AGEMA_reg_buffer_8982 ( .C (clk), .D (new_AGEMA_signal_21705), .Q (new_AGEMA_signal_21706) ) ;
    buf_clk new_AGEMA_reg_buffer_8985 ( .C (clk), .D (new_AGEMA_signal_21708), .Q (new_AGEMA_signal_21709) ) ;
    buf_clk new_AGEMA_reg_buffer_8988 ( .C (clk), .D (new_AGEMA_signal_21711), .Q (new_AGEMA_signal_21712) ) ;
    buf_clk new_AGEMA_reg_buffer_8991 ( .C (clk), .D (new_AGEMA_signal_21714), .Q (new_AGEMA_signal_21715) ) ;
    buf_clk new_AGEMA_reg_buffer_8994 ( .C (clk), .D (new_AGEMA_signal_21717), .Q (new_AGEMA_signal_21718) ) ;
    buf_clk new_AGEMA_reg_buffer_8997 ( .C (clk), .D (new_AGEMA_signal_21720), .Q (new_AGEMA_signal_21721) ) ;
    buf_clk new_AGEMA_reg_buffer_9000 ( .C (clk), .D (new_AGEMA_signal_21723), .Q (new_AGEMA_signal_21724) ) ;
    buf_clk new_AGEMA_reg_buffer_9003 ( .C (clk), .D (new_AGEMA_signal_21726), .Q (new_AGEMA_signal_21727) ) ;
    buf_clk new_AGEMA_reg_buffer_9006 ( .C (clk), .D (new_AGEMA_signal_21729), .Q (new_AGEMA_signal_21730) ) ;
    buf_clk new_AGEMA_reg_buffer_9009 ( .C (clk), .D (new_AGEMA_signal_21732), .Q (new_AGEMA_signal_21733) ) ;
    buf_clk new_AGEMA_reg_buffer_9012 ( .C (clk), .D (new_AGEMA_signal_21735), .Q (new_AGEMA_signal_21736) ) ;
    buf_clk new_AGEMA_reg_buffer_9015 ( .C (clk), .D (new_AGEMA_signal_21738), .Q (new_AGEMA_signal_21739) ) ;
    buf_clk new_AGEMA_reg_buffer_9018 ( .C (clk), .D (new_AGEMA_signal_21741), .Q (new_AGEMA_signal_21742) ) ;
    buf_clk new_AGEMA_reg_buffer_9021 ( .C (clk), .D (new_AGEMA_signal_21744), .Q (new_AGEMA_signal_21745) ) ;
    buf_clk new_AGEMA_reg_buffer_9024 ( .C (clk), .D (new_AGEMA_signal_21747), .Q (new_AGEMA_signal_21748) ) ;
    buf_clk new_AGEMA_reg_buffer_9027 ( .C (clk), .D (new_AGEMA_signal_21750), .Q (new_AGEMA_signal_21751) ) ;
    buf_clk new_AGEMA_reg_buffer_9030 ( .C (clk), .D (new_AGEMA_signal_21753), .Q (new_AGEMA_signal_21754) ) ;
    buf_clk new_AGEMA_reg_buffer_9033 ( .C (clk), .D (new_AGEMA_signal_21756), .Q (new_AGEMA_signal_21757) ) ;
    buf_clk new_AGEMA_reg_buffer_9036 ( .C (clk), .D (new_AGEMA_signal_21759), .Q (new_AGEMA_signal_21760) ) ;
    buf_clk new_AGEMA_reg_buffer_9039 ( .C (clk), .D (new_AGEMA_signal_21762), .Q (new_AGEMA_signal_21763) ) ;
    buf_clk new_AGEMA_reg_buffer_9042 ( .C (clk), .D (new_AGEMA_signal_21765), .Q (new_AGEMA_signal_21766) ) ;
    buf_clk new_AGEMA_reg_buffer_9045 ( .C (clk), .D (new_AGEMA_signal_21768), .Q (new_AGEMA_signal_21769) ) ;
    buf_clk new_AGEMA_reg_buffer_9048 ( .C (clk), .D (new_AGEMA_signal_21771), .Q (new_AGEMA_signal_21772) ) ;
    buf_clk new_AGEMA_reg_buffer_9051 ( .C (clk), .D (new_AGEMA_signal_21774), .Q (new_AGEMA_signal_21775) ) ;
    buf_clk new_AGEMA_reg_buffer_9054 ( .C (clk), .D (new_AGEMA_signal_21777), .Q (new_AGEMA_signal_21778) ) ;
    buf_clk new_AGEMA_reg_buffer_9057 ( .C (clk), .D (new_AGEMA_signal_21780), .Q (new_AGEMA_signal_21781) ) ;
    buf_clk new_AGEMA_reg_buffer_9060 ( .C (clk), .D (new_AGEMA_signal_21783), .Q (new_AGEMA_signal_21784) ) ;
    buf_clk new_AGEMA_reg_buffer_9063 ( .C (clk), .D (new_AGEMA_signal_21786), .Q (new_AGEMA_signal_21787) ) ;
    buf_clk new_AGEMA_reg_buffer_9066 ( .C (clk), .D (new_AGEMA_signal_21789), .Q (new_AGEMA_signal_21790) ) ;
    buf_clk new_AGEMA_reg_buffer_9069 ( .C (clk), .D (new_AGEMA_signal_21792), .Q (new_AGEMA_signal_21793) ) ;
    buf_clk new_AGEMA_reg_buffer_9072 ( .C (clk), .D (new_AGEMA_signal_21795), .Q (new_AGEMA_signal_21796) ) ;
    buf_clk new_AGEMA_reg_buffer_9075 ( .C (clk), .D (new_AGEMA_signal_21798), .Q (new_AGEMA_signal_21799) ) ;
    buf_clk new_AGEMA_reg_buffer_9078 ( .C (clk), .D (new_AGEMA_signal_21801), .Q (new_AGEMA_signal_21802) ) ;
    buf_clk new_AGEMA_reg_buffer_9081 ( .C (clk), .D (new_AGEMA_signal_21804), .Q (new_AGEMA_signal_21805) ) ;
    buf_clk new_AGEMA_reg_buffer_9084 ( .C (clk), .D (new_AGEMA_signal_21807), .Q (new_AGEMA_signal_21808) ) ;
    buf_clk new_AGEMA_reg_buffer_9087 ( .C (clk), .D (new_AGEMA_signal_21810), .Q (new_AGEMA_signal_21811) ) ;
    buf_clk new_AGEMA_reg_buffer_9090 ( .C (clk), .D (new_AGEMA_signal_21813), .Q (new_AGEMA_signal_21814) ) ;
    buf_clk new_AGEMA_reg_buffer_9094 ( .C (clk), .D (new_AGEMA_signal_21817), .Q (new_AGEMA_signal_21818) ) ;
    buf_clk new_AGEMA_reg_buffer_9098 ( .C (clk), .D (new_AGEMA_signal_21821), .Q (new_AGEMA_signal_21822) ) ;
    buf_clk new_AGEMA_reg_buffer_9102 ( .C (clk), .D (new_AGEMA_signal_21825), .Q (new_AGEMA_signal_21826) ) ;
    buf_clk new_AGEMA_reg_buffer_9106 ( .C (clk), .D (new_AGEMA_signal_21829), .Q (new_AGEMA_signal_21830) ) ;
    buf_clk new_AGEMA_reg_buffer_9110 ( .C (clk), .D (new_AGEMA_signal_21833), .Q (new_AGEMA_signal_21834) ) ;
    buf_clk new_AGEMA_reg_buffer_9114 ( .C (clk), .D (new_AGEMA_signal_21837), .Q (new_AGEMA_signal_21838) ) ;
    buf_clk new_AGEMA_reg_buffer_9118 ( .C (clk), .D (new_AGEMA_signal_21841), .Q (new_AGEMA_signal_21842) ) ;
    buf_clk new_AGEMA_reg_buffer_9122 ( .C (clk), .D (new_AGEMA_signal_21845), .Q (new_AGEMA_signal_21846) ) ;
    buf_clk new_AGEMA_reg_buffer_9126 ( .C (clk), .D (new_AGEMA_signal_21849), .Q (new_AGEMA_signal_21850) ) ;
    buf_clk new_AGEMA_reg_buffer_9130 ( .C (clk), .D (new_AGEMA_signal_21853), .Q (new_AGEMA_signal_21854) ) ;
    buf_clk new_AGEMA_reg_buffer_9134 ( .C (clk), .D (new_AGEMA_signal_21857), .Q (new_AGEMA_signal_21858) ) ;
    buf_clk new_AGEMA_reg_buffer_9138 ( .C (clk), .D (new_AGEMA_signal_21861), .Q (new_AGEMA_signal_21862) ) ;
    buf_clk new_AGEMA_reg_buffer_9142 ( .C (clk), .D (new_AGEMA_signal_21865), .Q (new_AGEMA_signal_21866) ) ;
    buf_clk new_AGEMA_reg_buffer_9146 ( .C (clk), .D (new_AGEMA_signal_21869), .Q (new_AGEMA_signal_21870) ) ;
    buf_clk new_AGEMA_reg_buffer_9150 ( .C (clk), .D (new_AGEMA_signal_21873), .Q (new_AGEMA_signal_21874) ) ;
    buf_clk new_AGEMA_reg_buffer_9154 ( .C (clk), .D (new_AGEMA_signal_21877), .Q (new_AGEMA_signal_21878) ) ;
    buf_clk new_AGEMA_reg_buffer_9158 ( .C (clk), .D (new_AGEMA_signal_21881), .Q (new_AGEMA_signal_21882) ) ;
    buf_clk new_AGEMA_reg_buffer_9162 ( .C (clk), .D (new_AGEMA_signal_21885), .Q (new_AGEMA_signal_21886) ) ;
    buf_clk new_AGEMA_reg_buffer_9166 ( .C (clk), .D (new_AGEMA_signal_21889), .Q (new_AGEMA_signal_21890) ) ;
    buf_clk new_AGEMA_reg_buffer_9170 ( .C (clk), .D (new_AGEMA_signal_21893), .Q (new_AGEMA_signal_21894) ) ;
    buf_clk new_AGEMA_reg_buffer_9174 ( .C (clk), .D (new_AGEMA_signal_21897), .Q (new_AGEMA_signal_21898) ) ;
    buf_clk new_AGEMA_reg_buffer_9178 ( .C (clk), .D (new_AGEMA_signal_21901), .Q (new_AGEMA_signal_21902) ) ;
    buf_clk new_AGEMA_reg_buffer_9182 ( .C (clk), .D (new_AGEMA_signal_21905), .Q (new_AGEMA_signal_21906) ) ;
    buf_clk new_AGEMA_reg_buffer_9186 ( .C (clk), .D (new_AGEMA_signal_21909), .Q (new_AGEMA_signal_21910) ) ;
    buf_clk new_AGEMA_reg_buffer_9190 ( .C (clk), .D (new_AGEMA_signal_21913), .Q (new_AGEMA_signal_21914) ) ;
    buf_clk new_AGEMA_reg_buffer_9194 ( .C (clk), .D (new_AGEMA_signal_21917), .Q (new_AGEMA_signal_21918) ) ;
    buf_clk new_AGEMA_reg_buffer_9198 ( .C (clk), .D (new_AGEMA_signal_21921), .Q (new_AGEMA_signal_21922) ) ;
    buf_clk new_AGEMA_reg_buffer_9202 ( .C (clk), .D (new_AGEMA_signal_21925), .Q (new_AGEMA_signal_21926) ) ;
    buf_clk new_AGEMA_reg_buffer_9206 ( .C (clk), .D (new_AGEMA_signal_21929), .Q (new_AGEMA_signal_21930) ) ;
    buf_clk new_AGEMA_reg_buffer_9210 ( .C (clk), .D (new_AGEMA_signal_21933), .Q (new_AGEMA_signal_21934) ) ;
    buf_clk new_AGEMA_reg_buffer_9214 ( .C (clk), .D (new_AGEMA_signal_21937), .Q (new_AGEMA_signal_21938) ) ;
    buf_clk new_AGEMA_reg_buffer_9218 ( .C (clk), .D (new_AGEMA_signal_21941), .Q (new_AGEMA_signal_21942) ) ;
    buf_clk new_AGEMA_reg_buffer_9222 ( .C (clk), .D (new_AGEMA_signal_21945), .Q (new_AGEMA_signal_21946) ) ;
    buf_clk new_AGEMA_reg_buffer_9226 ( .C (clk), .D (new_AGEMA_signal_21949), .Q (new_AGEMA_signal_21950) ) ;
    buf_clk new_AGEMA_reg_buffer_9230 ( .C (clk), .D (new_AGEMA_signal_21953), .Q (new_AGEMA_signal_21954) ) ;
    buf_clk new_AGEMA_reg_buffer_9234 ( .C (clk), .D (new_AGEMA_signal_21957), .Q (new_AGEMA_signal_21958) ) ;
    buf_clk new_AGEMA_reg_buffer_9238 ( .C (clk), .D (new_AGEMA_signal_21961), .Q (new_AGEMA_signal_21962) ) ;
    buf_clk new_AGEMA_reg_buffer_9242 ( .C (clk), .D (new_AGEMA_signal_21965), .Q (new_AGEMA_signal_21966) ) ;
    buf_clk new_AGEMA_reg_buffer_9246 ( .C (clk), .D (new_AGEMA_signal_21969), .Q (new_AGEMA_signal_21970) ) ;
    buf_clk new_AGEMA_reg_buffer_9250 ( .C (clk), .D (new_AGEMA_signal_21973), .Q (new_AGEMA_signal_21974) ) ;
    buf_clk new_AGEMA_reg_buffer_9254 ( .C (clk), .D (new_AGEMA_signal_21977), .Q (new_AGEMA_signal_21978) ) ;
    buf_clk new_AGEMA_reg_buffer_9258 ( .C (clk), .D (new_AGEMA_signal_21981), .Q (new_AGEMA_signal_21982) ) ;
    buf_clk new_AGEMA_reg_buffer_9262 ( .C (clk), .D (new_AGEMA_signal_21985), .Q (new_AGEMA_signal_21986) ) ;
    buf_clk new_AGEMA_reg_buffer_9266 ( .C (clk), .D (new_AGEMA_signal_21989), .Q (new_AGEMA_signal_21990) ) ;
    buf_clk new_AGEMA_reg_buffer_9270 ( .C (clk), .D (new_AGEMA_signal_21993), .Q (new_AGEMA_signal_21994) ) ;
    buf_clk new_AGEMA_reg_buffer_9274 ( .C (clk), .D (new_AGEMA_signal_21997), .Q (new_AGEMA_signal_21998) ) ;
    buf_clk new_AGEMA_reg_buffer_9278 ( .C (clk), .D (new_AGEMA_signal_22001), .Q (new_AGEMA_signal_22002) ) ;
    buf_clk new_AGEMA_reg_buffer_9282 ( .C (clk), .D (new_AGEMA_signal_22005), .Q (new_AGEMA_signal_22006) ) ;
    buf_clk new_AGEMA_reg_buffer_9286 ( .C (clk), .D (new_AGEMA_signal_22009), .Q (new_AGEMA_signal_22010) ) ;
    buf_clk new_AGEMA_reg_buffer_9290 ( .C (clk), .D (new_AGEMA_signal_22013), .Q (new_AGEMA_signal_22014) ) ;
    buf_clk new_AGEMA_reg_buffer_9294 ( .C (clk), .D (new_AGEMA_signal_22017), .Q (new_AGEMA_signal_22018) ) ;
    buf_clk new_AGEMA_reg_buffer_9298 ( .C (clk), .D (new_AGEMA_signal_22021), .Q (new_AGEMA_signal_22022) ) ;
    buf_clk new_AGEMA_reg_buffer_9302 ( .C (clk), .D (new_AGEMA_signal_22025), .Q (new_AGEMA_signal_22026) ) ;
    buf_clk new_AGEMA_reg_buffer_9306 ( .C (clk), .D (new_AGEMA_signal_22029), .Q (new_AGEMA_signal_22030) ) ;
    buf_clk new_AGEMA_reg_buffer_9310 ( .C (clk), .D (new_AGEMA_signal_22033), .Q (new_AGEMA_signal_22034) ) ;
    buf_clk new_AGEMA_reg_buffer_9314 ( .C (clk), .D (new_AGEMA_signal_22037), .Q (new_AGEMA_signal_22038) ) ;
    buf_clk new_AGEMA_reg_buffer_9318 ( .C (clk), .D (new_AGEMA_signal_22041), .Q (new_AGEMA_signal_22042) ) ;
    buf_clk new_AGEMA_reg_buffer_9322 ( .C (clk), .D (new_AGEMA_signal_22045), .Q (new_AGEMA_signal_22046) ) ;
    buf_clk new_AGEMA_reg_buffer_9326 ( .C (clk), .D (new_AGEMA_signal_22049), .Q (new_AGEMA_signal_22050) ) ;
    buf_clk new_AGEMA_reg_buffer_9330 ( .C (clk), .D (new_AGEMA_signal_22053), .Q (new_AGEMA_signal_22054) ) ;
    buf_clk new_AGEMA_reg_buffer_9334 ( .C (clk), .D (new_AGEMA_signal_22057), .Q (new_AGEMA_signal_22058) ) ;
    buf_clk new_AGEMA_reg_buffer_9338 ( .C (clk), .D (new_AGEMA_signal_22061), .Q (new_AGEMA_signal_22062) ) ;
    buf_clk new_AGEMA_reg_buffer_9342 ( .C (clk), .D (new_AGEMA_signal_22065), .Q (new_AGEMA_signal_22066) ) ;
    buf_clk new_AGEMA_reg_buffer_9346 ( .C (clk), .D (new_AGEMA_signal_22069), .Q (new_AGEMA_signal_22070) ) ;
    buf_clk new_AGEMA_reg_buffer_9350 ( .C (clk), .D (new_AGEMA_signal_22073), .Q (new_AGEMA_signal_22074) ) ;
    buf_clk new_AGEMA_reg_buffer_9354 ( .C (clk), .D (new_AGEMA_signal_22077), .Q (new_AGEMA_signal_22078) ) ;
    buf_clk new_AGEMA_reg_buffer_9358 ( .C (clk), .D (new_AGEMA_signal_22081), .Q (new_AGEMA_signal_22082) ) ;
    buf_clk new_AGEMA_reg_buffer_9362 ( .C (clk), .D (new_AGEMA_signal_22085), .Q (new_AGEMA_signal_22086) ) ;
    buf_clk new_AGEMA_reg_buffer_9366 ( .C (clk), .D (new_AGEMA_signal_22089), .Q (new_AGEMA_signal_22090) ) ;
    buf_clk new_AGEMA_reg_buffer_9370 ( .C (clk), .D (new_AGEMA_signal_22093), .Q (new_AGEMA_signal_22094) ) ;
    buf_clk new_AGEMA_reg_buffer_9374 ( .C (clk), .D (new_AGEMA_signal_22097), .Q (new_AGEMA_signal_22098) ) ;
    buf_clk new_AGEMA_reg_buffer_9378 ( .C (clk), .D (new_AGEMA_signal_22101), .Q (new_AGEMA_signal_22102) ) ;
    buf_clk new_AGEMA_reg_buffer_9382 ( .C (clk), .D (new_AGEMA_signal_22105), .Q (new_AGEMA_signal_22106) ) ;
    buf_clk new_AGEMA_reg_buffer_9386 ( .C (clk), .D (new_AGEMA_signal_22109), .Q (new_AGEMA_signal_22110) ) ;
    buf_clk new_AGEMA_reg_buffer_9390 ( .C (clk), .D (new_AGEMA_signal_22113), .Q (new_AGEMA_signal_22114) ) ;
    buf_clk new_AGEMA_reg_buffer_9394 ( .C (clk), .D (new_AGEMA_signal_22117), .Q (new_AGEMA_signal_22118) ) ;
    buf_clk new_AGEMA_reg_buffer_9398 ( .C (clk), .D (new_AGEMA_signal_22121), .Q (new_AGEMA_signal_22122) ) ;
    buf_clk new_AGEMA_reg_buffer_9402 ( .C (clk), .D (new_AGEMA_signal_22125), .Q (new_AGEMA_signal_22126) ) ;
    buf_clk new_AGEMA_reg_buffer_9406 ( .C (clk), .D (new_AGEMA_signal_22129), .Q (new_AGEMA_signal_22130) ) ;
    buf_clk new_AGEMA_reg_buffer_9410 ( .C (clk), .D (new_AGEMA_signal_22133), .Q (new_AGEMA_signal_22134) ) ;
    buf_clk new_AGEMA_reg_buffer_9414 ( .C (clk), .D (new_AGEMA_signal_22137), .Q (new_AGEMA_signal_22138) ) ;
    buf_clk new_AGEMA_reg_buffer_9418 ( .C (clk), .D (new_AGEMA_signal_22141), .Q (new_AGEMA_signal_22142) ) ;
    buf_clk new_AGEMA_reg_buffer_9422 ( .C (clk), .D (new_AGEMA_signal_22145), .Q (new_AGEMA_signal_22146) ) ;
    buf_clk new_AGEMA_reg_buffer_9426 ( .C (clk), .D (new_AGEMA_signal_22149), .Q (new_AGEMA_signal_22150) ) ;
    buf_clk new_AGEMA_reg_buffer_9430 ( .C (clk), .D (new_AGEMA_signal_22153), .Q (new_AGEMA_signal_22154) ) ;
    buf_clk new_AGEMA_reg_buffer_9434 ( .C (clk), .D (new_AGEMA_signal_22157), .Q (new_AGEMA_signal_22158) ) ;
    buf_clk new_AGEMA_reg_buffer_9438 ( .C (clk), .D (new_AGEMA_signal_22161), .Q (new_AGEMA_signal_22162) ) ;
    buf_clk new_AGEMA_reg_buffer_9442 ( .C (clk), .D (new_AGEMA_signal_22165), .Q (new_AGEMA_signal_22166) ) ;
    buf_clk new_AGEMA_reg_buffer_9446 ( .C (clk), .D (new_AGEMA_signal_22169), .Q (new_AGEMA_signal_22170) ) ;
    buf_clk new_AGEMA_reg_buffer_9450 ( .C (clk), .D (new_AGEMA_signal_22173), .Q (new_AGEMA_signal_22174) ) ;
    buf_clk new_AGEMA_reg_buffer_9454 ( .C (clk), .D (new_AGEMA_signal_22177), .Q (new_AGEMA_signal_22178) ) ;
    buf_clk new_AGEMA_reg_buffer_9458 ( .C (clk), .D (new_AGEMA_signal_22181), .Q (new_AGEMA_signal_22182) ) ;
    buf_clk new_AGEMA_reg_buffer_9462 ( .C (clk), .D (new_AGEMA_signal_22185), .Q (new_AGEMA_signal_22186) ) ;
    buf_clk new_AGEMA_reg_buffer_9466 ( .C (clk), .D (new_AGEMA_signal_22189), .Q (new_AGEMA_signal_22190) ) ;
    buf_clk new_AGEMA_reg_buffer_9470 ( .C (clk), .D (new_AGEMA_signal_22193), .Q (new_AGEMA_signal_22194) ) ;
    buf_clk new_AGEMA_reg_buffer_9474 ( .C (clk), .D (new_AGEMA_signal_22197), .Q (new_AGEMA_signal_22198) ) ;
    buf_clk new_AGEMA_reg_buffer_9478 ( .C (clk), .D (new_AGEMA_signal_22201), .Q (new_AGEMA_signal_22202) ) ;
    buf_clk new_AGEMA_reg_buffer_9482 ( .C (clk), .D (new_AGEMA_signal_22205), .Q (new_AGEMA_signal_22206) ) ;
    buf_clk new_AGEMA_reg_buffer_9486 ( .C (clk), .D (new_AGEMA_signal_22209), .Q (new_AGEMA_signal_22210) ) ;
    buf_clk new_AGEMA_reg_buffer_9490 ( .C (clk), .D (new_AGEMA_signal_22213), .Q (new_AGEMA_signal_22214) ) ;
    buf_clk new_AGEMA_reg_buffer_9494 ( .C (clk), .D (new_AGEMA_signal_22217), .Q (new_AGEMA_signal_22218) ) ;
    buf_clk new_AGEMA_reg_buffer_9498 ( .C (clk), .D (new_AGEMA_signal_22221), .Q (new_AGEMA_signal_22222) ) ;
    buf_clk new_AGEMA_reg_buffer_9502 ( .C (clk), .D (new_AGEMA_signal_22225), .Q (new_AGEMA_signal_22226) ) ;
    buf_clk new_AGEMA_reg_buffer_9506 ( .C (clk), .D (new_AGEMA_signal_22229), .Q (new_AGEMA_signal_22230) ) ;
    buf_clk new_AGEMA_reg_buffer_9510 ( .C (clk), .D (new_AGEMA_signal_22233), .Q (new_AGEMA_signal_22234) ) ;
    buf_clk new_AGEMA_reg_buffer_9514 ( .C (clk), .D (new_AGEMA_signal_22237), .Q (new_AGEMA_signal_22238) ) ;
    buf_clk new_AGEMA_reg_buffer_9518 ( .C (clk), .D (new_AGEMA_signal_22241), .Q (new_AGEMA_signal_22242) ) ;
    buf_clk new_AGEMA_reg_buffer_9522 ( .C (clk), .D (new_AGEMA_signal_22245), .Q (new_AGEMA_signal_22246) ) ;
    buf_clk new_AGEMA_reg_buffer_9526 ( .C (clk), .D (new_AGEMA_signal_22249), .Q (new_AGEMA_signal_22250) ) ;
    buf_clk new_AGEMA_reg_buffer_9530 ( .C (clk), .D (new_AGEMA_signal_22253), .Q (new_AGEMA_signal_22254) ) ;
    buf_clk new_AGEMA_reg_buffer_9534 ( .C (clk), .D (new_AGEMA_signal_22257), .Q (new_AGEMA_signal_22258) ) ;
    buf_clk new_AGEMA_reg_buffer_9538 ( .C (clk), .D (new_AGEMA_signal_22261), .Q (new_AGEMA_signal_22262) ) ;
    buf_clk new_AGEMA_reg_buffer_9542 ( .C (clk), .D (new_AGEMA_signal_22265), .Q (new_AGEMA_signal_22266) ) ;
    buf_clk new_AGEMA_reg_buffer_9546 ( .C (clk), .D (new_AGEMA_signal_22269), .Q (new_AGEMA_signal_22270) ) ;
    buf_clk new_AGEMA_reg_buffer_9550 ( .C (clk), .D (new_AGEMA_signal_22273), .Q (new_AGEMA_signal_22274) ) ;
    buf_clk new_AGEMA_reg_buffer_9554 ( .C (clk), .D (new_AGEMA_signal_22277), .Q (new_AGEMA_signal_22278) ) ;
    buf_clk new_AGEMA_reg_buffer_9558 ( .C (clk), .D (new_AGEMA_signal_22281), .Q (new_AGEMA_signal_22282) ) ;
    buf_clk new_AGEMA_reg_buffer_9562 ( .C (clk), .D (new_AGEMA_signal_22285), .Q (new_AGEMA_signal_22286) ) ;
    buf_clk new_AGEMA_reg_buffer_9566 ( .C (clk), .D (new_AGEMA_signal_22289), .Q (new_AGEMA_signal_22290) ) ;
    buf_clk new_AGEMA_reg_buffer_9570 ( .C (clk), .D (new_AGEMA_signal_22293), .Q (new_AGEMA_signal_22294) ) ;
    buf_clk new_AGEMA_reg_buffer_9574 ( .C (clk), .D (new_AGEMA_signal_22297), .Q (new_AGEMA_signal_22298) ) ;
    buf_clk new_AGEMA_reg_buffer_9578 ( .C (clk), .D (new_AGEMA_signal_22301), .Q (new_AGEMA_signal_22302) ) ;
    buf_clk new_AGEMA_reg_buffer_9582 ( .C (clk), .D (new_AGEMA_signal_22305), .Q (new_AGEMA_signal_22306) ) ;
    buf_clk new_AGEMA_reg_buffer_9586 ( .C (clk), .D (new_AGEMA_signal_22309), .Q (new_AGEMA_signal_22310) ) ;
    buf_clk new_AGEMA_reg_buffer_9590 ( .C (clk), .D (new_AGEMA_signal_22313), .Q (new_AGEMA_signal_22314) ) ;
    buf_clk new_AGEMA_reg_buffer_9594 ( .C (clk), .D (new_AGEMA_signal_22317), .Q (new_AGEMA_signal_22318) ) ;
    buf_clk new_AGEMA_reg_buffer_9598 ( .C (clk), .D (new_AGEMA_signal_22321), .Q (new_AGEMA_signal_22322) ) ;
    buf_clk new_AGEMA_reg_buffer_9602 ( .C (clk), .D (new_AGEMA_signal_22325), .Q (new_AGEMA_signal_22326) ) ;
    buf_clk new_AGEMA_reg_buffer_9606 ( .C (clk), .D (new_AGEMA_signal_22329), .Q (new_AGEMA_signal_22330) ) ;
    buf_clk new_AGEMA_reg_buffer_9610 ( .C (clk), .D (new_AGEMA_signal_22333), .Q (new_AGEMA_signal_22334) ) ;
    buf_clk new_AGEMA_reg_buffer_9614 ( .C (clk), .D (new_AGEMA_signal_22337), .Q (new_AGEMA_signal_22338) ) ;
    buf_clk new_AGEMA_reg_buffer_9618 ( .C (clk), .D (new_AGEMA_signal_22341), .Q (new_AGEMA_signal_22342) ) ;
    buf_clk new_AGEMA_reg_buffer_9622 ( .C (clk), .D (new_AGEMA_signal_22345), .Q (new_AGEMA_signal_22346) ) ;
    buf_clk new_AGEMA_reg_buffer_9626 ( .C (clk), .D (new_AGEMA_signal_22349), .Q (new_AGEMA_signal_22350) ) ;
    buf_clk new_AGEMA_reg_buffer_9630 ( .C (clk), .D (new_AGEMA_signal_22353), .Q (new_AGEMA_signal_22354) ) ;
    buf_clk new_AGEMA_reg_buffer_9634 ( .C (clk), .D (new_AGEMA_signal_22357), .Q (new_AGEMA_signal_22358) ) ;
    buf_clk new_AGEMA_reg_buffer_9638 ( .C (clk), .D (new_AGEMA_signal_22361), .Q (new_AGEMA_signal_22362) ) ;
    buf_clk new_AGEMA_reg_buffer_9642 ( .C (clk), .D (new_AGEMA_signal_22365), .Q (new_AGEMA_signal_22366) ) ;
    buf_clk new_AGEMA_reg_buffer_9646 ( .C (clk), .D (new_AGEMA_signal_22369), .Q (new_AGEMA_signal_22370) ) ;
    buf_clk new_AGEMA_reg_buffer_9650 ( .C (clk), .D (new_AGEMA_signal_22373), .Q (new_AGEMA_signal_22374) ) ;
    buf_clk new_AGEMA_reg_buffer_9654 ( .C (clk), .D (new_AGEMA_signal_22377), .Q (new_AGEMA_signal_22378) ) ;
    buf_clk new_AGEMA_reg_buffer_9658 ( .C (clk), .D (new_AGEMA_signal_22381), .Q (new_AGEMA_signal_22382) ) ;
    buf_clk new_AGEMA_reg_buffer_9662 ( .C (clk), .D (new_AGEMA_signal_22385), .Q (new_AGEMA_signal_22386) ) ;
    buf_clk new_AGEMA_reg_buffer_9666 ( .C (clk), .D (new_AGEMA_signal_22389), .Q (new_AGEMA_signal_22390) ) ;
    buf_clk new_AGEMA_reg_buffer_9670 ( .C (clk), .D (new_AGEMA_signal_22393), .Q (new_AGEMA_signal_22394) ) ;
    buf_clk new_AGEMA_reg_buffer_9674 ( .C (clk), .D (new_AGEMA_signal_22397), .Q (new_AGEMA_signal_22398) ) ;
    buf_clk new_AGEMA_reg_buffer_9678 ( .C (clk), .D (new_AGEMA_signal_22401), .Q (new_AGEMA_signal_22402) ) ;
    buf_clk new_AGEMA_reg_buffer_9682 ( .C (clk), .D (new_AGEMA_signal_22405), .Q (new_AGEMA_signal_22406) ) ;
    buf_clk new_AGEMA_reg_buffer_9686 ( .C (clk), .D (new_AGEMA_signal_22409), .Q (new_AGEMA_signal_22410) ) ;
    buf_clk new_AGEMA_reg_buffer_9690 ( .C (clk), .D (new_AGEMA_signal_22413), .Q (new_AGEMA_signal_22414) ) ;
    buf_clk new_AGEMA_reg_buffer_9694 ( .C (clk), .D (new_AGEMA_signal_22417), .Q (new_AGEMA_signal_22418) ) ;
    buf_clk new_AGEMA_reg_buffer_9698 ( .C (clk), .D (new_AGEMA_signal_22421), .Q (new_AGEMA_signal_22422) ) ;
    buf_clk new_AGEMA_reg_buffer_9702 ( .C (clk), .D (new_AGEMA_signal_22425), .Q (new_AGEMA_signal_22426) ) ;
    buf_clk new_AGEMA_reg_buffer_9706 ( .C (clk), .D (new_AGEMA_signal_22429), .Q (new_AGEMA_signal_22430) ) ;
    buf_clk new_AGEMA_reg_buffer_9710 ( .C (clk), .D (new_AGEMA_signal_22433), .Q (new_AGEMA_signal_22434) ) ;
    buf_clk new_AGEMA_reg_buffer_9714 ( .C (clk), .D (new_AGEMA_signal_22437), .Q (new_AGEMA_signal_22438) ) ;
    buf_clk new_AGEMA_reg_buffer_9718 ( .C (clk), .D (new_AGEMA_signal_22441), .Q (new_AGEMA_signal_22442) ) ;
    buf_clk new_AGEMA_reg_buffer_9722 ( .C (clk), .D (new_AGEMA_signal_22445), .Q (new_AGEMA_signal_22446) ) ;
    buf_clk new_AGEMA_reg_buffer_9726 ( .C (clk), .D (new_AGEMA_signal_22449), .Q (new_AGEMA_signal_22450) ) ;
    buf_clk new_AGEMA_reg_buffer_9730 ( .C (clk), .D (new_AGEMA_signal_22453), .Q (new_AGEMA_signal_22454) ) ;
    buf_clk new_AGEMA_reg_buffer_9734 ( .C (clk), .D (new_AGEMA_signal_22457), .Q (new_AGEMA_signal_22458) ) ;
    buf_clk new_AGEMA_reg_buffer_9738 ( .C (clk), .D (new_AGEMA_signal_22461), .Q (new_AGEMA_signal_22462) ) ;
    buf_clk new_AGEMA_reg_buffer_9742 ( .C (clk), .D (new_AGEMA_signal_22465), .Q (new_AGEMA_signal_22466) ) ;
    buf_clk new_AGEMA_reg_buffer_9746 ( .C (clk), .D (new_AGEMA_signal_22469), .Q (new_AGEMA_signal_22470) ) ;
    buf_clk new_AGEMA_reg_buffer_9750 ( .C (clk), .D (new_AGEMA_signal_22473), .Q (new_AGEMA_signal_22474) ) ;
    buf_clk new_AGEMA_reg_buffer_9754 ( .C (clk), .D (new_AGEMA_signal_22477), .Q (new_AGEMA_signal_22478) ) ;
    buf_clk new_AGEMA_reg_buffer_9758 ( .C (clk), .D (new_AGEMA_signal_22481), .Q (new_AGEMA_signal_22482) ) ;
    buf_clk new_AGEMA_reg_buffer_9762 ( .C (clk), .D (new_AGEMA_signal_22485), .Q (new_AGEMA_signal_22486) ) ;
    buf_clk new_AGEMA_reg_buffer_9766 ( .C (clk), .D (new_AGEMA_signal_22489), .Q (new_AGEMA_signal_22490) ) ;
    buf_clk new_AGEMA_reg_buffer_9770 ( .C (clk), .D (new_AGEMA_signal_22493), .Q (new_AGEMA_signal_22494) ) ;
    buf_clk new_AGEMA_reg_buffer_9774 ( .C (clk), .D (new_AGEMA_signal_22497), .Q (new_AGEMA_signal_22498) ) ;
    buf_clk new_AGEMA_reg_buffer_9778 ( .C (clk), .D (new_AGEMA_signal_22501), .Q (new_AGEMA_signal_22502) ) ;
    buf_clk new_AGEMA_reg_buffer_9782 ( .C (clk), .D (new_AGEMA_signal_22505), .Q (new_AGEMA_signal_22506) ) ;
    buf_clk new_AGEMA_reg_buffer_9786 ( .C (clk), .D (new_AGEMA_signal_22509), .Q (new_AGEMA_signal_22510) ) ;
    buf_clk new_AGEMA_reg_buffer_9790 ( .C (clk), .D (new_AGEMA_signal_22513), .Q (new_AGEMA_signal_22514) ) ;
    buf_clk new_AGEMA_reg_buffer_9794 ( .C (clk), .D (new_AGEMA_signal_22517), .Q (new_AGEMA_signal_22518) ) ;
    buf_clk new_AGEMA_reg_buffer_9798 ( .C (clk), .D (new_AGEMA_signal_22521), .Q (new_AGEMA_signal_22522) ) ;
    buf_clk new_AGEMA_reg_buffer_9802 ( .C (clk), .D (new_AGEMA_signal_22525), .Q (new_AGEMA_signal_22526) ) ;
    buf_clk new_AGEMA_reg_buffer_9806 ( .C (clk), .D (new_AGEMA_signal_22529), .Q (new_AGEMA_signal_22530) ) ;
    buf_clk new_AGEMA_reg_buffer_9810 ( .C (clk), .D (new_AGEMA_signal_22533), .Q (new_AGEMA_signal_22534) ) ;
    buf_clk new_AGEMA_reg_buffer_9814 ( .C (clk), .D (new_AGEMA_signal_22537), .Q (new_AGEMA_signal_22538) ) ;
    buf_clk new_AGEMA_reg_buffer_9818 ( .C (clk), .D (new_AGEMA_signal_22541), .Q (new_AGEMA_signal_22542) ) ;
    buf_clk new_AGEMA_reg_buffer_9822 ( .C (clk), .D (new_AGEMA_signal_22545), .Q (new_AGEMA_signal_22546) ) ;
    buf_clk new_AGEMA_reg_buffer_9826 ( .C (clk), .D (new_AGEMA_signal_22549), .Q (new_AGEMA_signal_22550) ) ;
    buf_clk new_AGEMA_reg_buffer_9830 ( .C (clk), .D (new_AGEMA_signal_22553), .Q (new_AGEMA_signal_22554) ) ;
    buf_clk new_AGEMA_reg_buffer_9834 ( .C (clk), .D (new_AGEMA_signal_22557), .Q (new_AGEMA_signal_22558) ) ;
    buf_clk new_AGEMA_reg_buffer_9838 ( .C (clk), .D (new_AGEMA_signal_22561), .Q (new_AGEMA_signal_22562) ) ;
    buf_clk new_AGEMA_reg_buffer_9842 ( .C (clk), .D (new_AGEMA_signal_22565), .Q (new_AGEMA_signal_22566) ) ;
    buf_clk new_AGEMA_reg_buffer_9846 ( .C (clk), .D (new_AGEMA_signal_22569), .Q (new_AGEMA_signal_22570) ) ;
    buf_clk new_AGEMA_reg_buffer_9850 ( .C (clk), .D (new_AGEMA_signal_22573), .Q (new_AGEMA_signal_22574) ) ;
    buf_clk new_AGEMA_reg_buffer_9854 ( .C (clk), .D (new_AGEMA_signal_22577), .Q (new_AGEMA_signal_22578) ) ;
    buf_clk new_AGEMA_reg_buffer_9858 ( .C (clk), .D (new_AGEMA_signal_22581), .Q (new_AGEMA_signal_22582) ) ;
    buf_clk new_AGEMA_reg_buffer_9862 ( .C (clk), .D (new_AGEMA_signal_22585), .Q (new_AGEMA_signal_22586) ) ;
    buf_clk new_AGEMA_reg_buffer_9866 ( .C (clk), .D (new_AGEMA_signal_22589), .Q (new_AGEMA_signal_22590) ) ;
    buf_clk new_AGEMA_reg_buffer_9870 ( .C (clk), .D (new_AGEMA_signal_22593), .Q (new_AGEMA_signal_22594) ) ;
    buf_clk new_AGEMA_reg_buffer_9874 ( .C (clk), .D (new_AGEMA_signal_22597), .Q (new_AGEMA_signal_22598) ) ;
    buf_clk new_AGEMA_reg_buffer_9878 ( .C (clk), .D (new_AGEMA_signal_22601), .Q (new_AGEMA_signal_22602) ) ;
    buf_clk new_AGEMA_reg_buffer_9882 ( .C (clk), .D (new_AGEMA_signal_22605), .Q (new_AGEMA_signal_22606) ) ;
    buf_clk new_AGEMA_reg_buffer_9886 ( .C (clk), .D (new_AGEMA_signal_22609), .Q (new_AGEMA_signal_22610) ) ;
    buf_clk new_AGEMA_reg_buffer_9890 ( .C (clk), .D (new_AGEMA_signal_22613), .Q (new_AGEMA_signal_22614) ) ;
    buf_clk new_AGEMA_reg_buffer_9894 ( .C (clk), .D (new_AGEMA_signal_22617), .Q (new_AGEMA_signal_22618) ) ;
    buf_clk new_AGEMA_reg_buffer_9898 ( .C (clk), .D (new_AGEMA_signal_22621), .Q (new_AGEMA_signal_22622) ) ;
    buf_clk new_AGEMA_reg_buffer_9902 ( .C (clk), .D (new_AGEMA_signal_22625), .Q (new_AGEMA_signal_22626) ) ;
    buf_clk new_AGEMA_reg_buffer_9906 ( .C (clk), .D (new_AGEMA_signal_22629), .Q (new_AGEMA_signal_22630) ) ;
    buf_clk new_AGEMA_reg_buffer_9910 ( .C (clk), .D (new_AGEMA_signal_22633), .Q (new_AGEMA_signal_22634) ) ;
    buf_clk new_AGEMA_reg_buffer_9914 ( .C (clk), .D (new_AGEMA_signal_22637), .Q (new_AGEMA_signal_22638) ) ;
    buf_clk new_AGEMA_reg_buffer_9918 ( .C (clk), .D (new_AGEMA_signal_22641), .Q (new_AGEMA_signal_22642) ) ;
    buf_clk new_AGEMA_reg_buffer_9922 ( .C (clk), .D (new_AGEMA_signal_22645), .Q (new_AGEMA_signal_22646) ) ;
    buf_clk new_AGEMA_reg_buffer_9926 ( .C (clk), .D (new_AGEMA_signal_22649), .Q (new_AGEMA_signal_22650) ) ;
    buf_clk new_AGEMA_reg_buffer_9930 ( .C (clk), .D (new_AGEMA_signal_22653), .Q (new_AGEMA_signal_22654) ) ;
    buf_clk new_AGEMA_reg_buffer_9934 ( .C (clk), .D (new_AGEMA_signal_22657), .Q (new_AGEMA_signal_22658) ) ;
    buf_clk new_AGEMA_reg_buffer_9938 ( .C (clk), .D (new_AGEMA_signal_22661), .Q (new_AGEMA_signal_22662) ) ;
    buf_clk new_AGEMA_reg_buffer_9942 ( .C (clk), .D (new_AGEMA_signal_22665), .Q (new_AGEMA_signal_22666) ) ;
    buf_clk new_AGEMA_reg_buffer_9946 ( .C (clk), .D (new_AGEMA_signal_22669), .Q (new_AGEMA_signal_22670) ) ;
    buf_clk new_AGEMA_reg_buffer_9950 ( .C (clk), .D (new_AGEMA_signal_22673), .Q (new_AGEMA_signal_22674) ) ;
    buf_clk new_AGEMA_reg_buffer_9954 ( .C (clk), .D (new_AGEMA_signal_22677), .Q (new_AGEMA_signal_22678) ) ;
    buf_clk new_AGEMA_reg_buffer_9958 ( .C (clk), .D (new_AGEMA_signal_22681), .Q (new_AGEMA_signal_22682) ) ;
    buf_clk new_AGEMA_reg_buffer_9962 ( .C (clk), .D (new_AGEMA_signal_22685), .Q (new_AGEMA_signal_22686) ) ;
    buf_clk new_AGEMA_reg_buffer_9966 ( .C (clk), .D (new_AGEMA_signal_22689), .Q (new_AGEMA_signal_22690) ) ;
    buf_clk new_AGEMA_reg_buffer_9970 ( .C (clk), .D (new_AGEMA_signal_22693), .Q (new_AGEMA_signal_22694) ) ;
    buf_clk new_AGEMA_reg_buffer_9974 ( .C (clk), .D (new_AGEMA_signal_22697), .Q (new_AGEMA_signal_22698) ) ;
    buf_clk new_AGEMA_reg_buffer_9978 ( .C (clk), .D (new_AGEMA_signal_22701), .Q (new_AGEMA_signal_22702) ) ;
    buf_clk new_AGEMA_reg_buffer_9982 ( .C (clk), .D (new_AGEMA_signal_22705), .Q (new_AGEMA_signal_22706) ) ;
    buf_clk new_AGEMA_reg_buffer_9986 ( .C (clk), .D (new_AGEMA_signal_22709), .Q (new_AGEMA_signal_22710) ) ;
    buf_clk new_AGEMA_reg_buffer_9990 ( .C (clk), .D (new_AGEMA_signal_22713), .Q (new_AGEMA_signal_22714) ) ;
    buf_clk new_AGEMA_reg_buffer_9994 ( .C (clk), .D (new_AGEMA_signal_22717), .Q (new_AGEMA_signal_22718) ) ;
    buf_clk new_AGEMA_reg_buffer_9998 ( .C (clk), .D (new_AGEMA_signal_22721), .Q (new_AGEMA_signal_22722) ) ;
    buf_clk new_AGEMA_reg_buffer_10002 ( .C (clk), .D (new_AGEMA_signal_22725), .Q (new_AGEMA_signal_22726) ) ;
    buf_clk new_AGEMA_reg_buffer_10006 ( .C (clk), .D (new_AGEMA_signal_22729), .Q (new_AGEMA_signal_22730) ) ;
    buf_clk new_AGEMA_reg_buffer_10010 ( .C (clk), .D (new_AGEMA_signal_22733), .Q (new_AGEMA_signal_22734) ) ;
    buf_clk new_AGEMA_reg_buffer_10014 ( .C (clk), .D (new_AGEMA_signal_22737), .Q (new_AGEMA_signal_22738) ) ;
    buf_clk new_AGEMA_reg_buffer_10018 ( .C (clk), .D (new_AGEMA_signal_22741), .Q (new_AGEMA_signal_22742) ) ;
    buf_clk new_AGEMA_reg_buffer_10022 ( .C (clk), .D (new_AGEMA_signal_22745), .Q (new_AGEMA_signal_22746) ) ;
    buf_clk new_AGEMA_reg_buffer_10026 ( .C (clk), .D (new_AGEMA_signal_22749), .Q (new_AGEMA_signal_22750) ) ;
    buf_clk new_AGEMA_reg_buffer_10030 ( .C (clk), .D (new_AGEMA_signal_22753), .Q (new_AGEMA_signal_22754) ) ;
    buf_clk new_AGEMA_reg_buffer_10034 ( .C (clk), .D (new_AGEMA_signal_22757), .Q (new_AGEMA_signal_22758) ) ;
    buf_clk new_AGEMA_reg_buffer_10038 ( .C (clk), .D (new_AGEMA_signal_22761), .Q (new_AGEMA_signal_22762) ) ;
    buf_clk new_AGEMA_reg_buffer_10042 ( .C (clk), .D (new_AGEMA_signal_22765), .Q (new_AGEMA_signal_22766) ) ;
    buf_clk new_AGEMA_reg_buffer_10046 ( .C (clk), .D (new_AGEMA_signal_22769), .Q (new_AGEMA_signal_22770) ) ;
    buf_clk new_AGEMA_reg_buffer_10050 ( .C (clk), .D (new_AGEMA_signal_22773), .Q (new_AGEMA_signal_22774) ) ;
    buf_clk new_AGEMA_reg_buffer_10054 ( .C (clk), .D (new_AGEMA_signal_22777), .Q (new_AGEMA_signal_22778) ) ;
    buf_clk new_AGEMA_reg_buffer_10058 ( .C (clk), .D (new_AGEMA_signal_22781), .Q (new_AGEMA_signal_22782) ) ;
    buf_clk new_AGEMA_reg_buffer_10062 ( .C (clk), .D (new_AGEMA_signal_22785), .Q (new_AGEMA_signal_22786) ) ;
    buf_clk new_AGEMA_reg_buffer_10066 ( .C (clk), .D (new_AGEMA_signal_22789), .Q (new_AGEMA_signal_22790) ) ;
    buf_clk new_AGEMA_reg_buffer_10070 ( .C (clk), .D (new_AGEMA_signal_22793), .Q (new_AGEMA_signal_22794) ) ;
    buf_clk new_AGEMA_reg_buffer_10074 ( .C (clk), .D (new_AGEMA_signal_22797), .Q (new_AGEMA_signal_22798) ) ;
    buf_clk new_AGEMA_reg_buffer_10078 ( .C (clk), .D (new_AGEMA_signal_22801), .Q (new_AGEMA_signal_22802) ) ;
    buf_clk new_AGEMA_reg_buffer_10082 ( .C (clk), .D (new_AGEMA_signal_22805), .Q (new_AGEMA_signal_22806) ) ;
    buf_clk new_AGEMA_reg_buffer_10086 ( .C (clk), .D (new_AGEMA_signal_22809), .Q (new_AGEMA_signal_22810) ) ;
    buf_clk new_AGEMA_reg_buffer_10090 ( .C (clk), .D (new_AGEMA_signal_22813), .Q (new_AGEMA_signal_22814) ) ;
    buf_clk new_AGEMA_reg_buffer_10094 ( .C (clk), .D (new_AGEMA_signal_22817), .Q (new_AGEMA_signal_22818) ) ;
    buf_clk new_AGEMA_reg_buffer_10098 ( .C (clk), .D (new_AGEMA_signal_22821), .Q (new_AGEMA_signal_22822) ) ;
    buf_clk new_AGEMA_reg_buffer_10102 ( .C (clk), .D (new_AGEMA_signal_22825), .Q (new_AGEMA_signal_22826) ) ;
    buf_clk new_AGEMA_reg_buffer_10106 ( .C (clk), .D (new_AGEMA_signal_22829), .Q (new_AGEMA_signal_22830) ) ;
    buf_clk new_AGEMA_reg_buffer_10110 ( .C (clk), .D (new_AGEMA_signal_22833), .Q (new_AGEMA_signal_22834) ) ;
    buf_clk new_AGEMA_reg_buffer_10114 ( .C (clk), .D (new_AGEMA_signal_22837), .Q (new_AGEMA_signal_22838) ) ;
    buf_clk new_AGEMA_reg_buffer_10118 ( .C (clk), .D (new_AGEMA_signal_22841), .Q (new_AGEMA_signal_22842) ) ;
    buf_clk new_AGEMA_reg_buffer_10122 ( .C (clk), .D (new_AGEMA_signal_22845), .Q (new_AGEMA_signal_22846) ) ;
    buf_clk new_AGEMA_reg_buffer_10126 ( .C (clk), .D (new_AGEMA_signal_22849), .Q (new_AGEMA_signal_22850) ) ;
    buf_clk new_AGEMA_reg_buffer_10130 ( .C (clk), .D (new_AGEMA_signal_22853), .Q (new_AGEMA_signal_22854) ) ;
    buf_clk new_AGEMA_reg_buffer_10134 ( .C (clk), .D (new_AGEMA_signal_22857), .Q (new_AGEMA_signal_22858) ) ;
    buf_clk new_AGEMA_reg_buffer_10138 ( .C (clk), .D (new_AGEMA_signal_22861), .Q (new_AGEMA_signal_22862) ) ;
    buf_clk new_AGEMA_reg_buffer_10142 ( .C (clk), .D (new_AGEMA_signal_22865), .Q (new_AGEMA_signal_22866) ) ;
    buf_clk new_AGEMA_reg_buffer_10146 ( .C (clk), .D (new_AGEMA_signal_22869), .Q (new_AGEMA_signal_22870) ) ;
    buf_clk new_AGEMA_reg_buffer_10150 ( .C (clk), .D (new_AGEMA_signal_22873), .Q (new_AGEMA_signal_22874) ) ;
    buf_clk new_AGEMA_reg_buffer_10154 ( .C (clk), .D (new_AGEMA_signal_22877), .Q (new_AGEMA_signal_22878) ) ;
    buf_clk new_AGEMA_reg_buffer_10158 ( .C (clk), .D (new_AGEMA_signal_22881), .Q (new_AGEMA_signal_22882) ) ;
    buf_clk new_AGEMA_reg_buffer_10162 ( .C (clk), .D (new_AGEMA_signal_22885), .Q (new_AGEMA_signal_22886) ) ;
    buf_clk new_AGEMA_reg_buffer_10166 ( .C (clk), .D (new_AGEMA_signal_22889), .Q (new_AGEMA_signal_22890) ) ;
    buf_clk new_AGEMA_reg_buffer_10170 ( .C (clk), .D (new_AGEMA_signal_22893), .Q (new_AGEMA_signal_22894) ) ;
    buf_clk new_AGEMA_reg_buffer_10174 ( .C (clk), .D (new_AGEMA_signal_22897), .Q (new_AGEMA_signal_22898) ) ;
    buf_clk new_AGEMA_reg_buffer_10178 ( .C (clk), .D (new_AGEMA_signal_22901), .Q (new_AGEMA_signal_22902) ) ;
    buf_clk new_AGEMA_reg_buffer_10182 ( .C (clk), .D (new_AGEMA_signal_22905), .Q (new_AGEMA_signal_22906) ) ;
    buf_clk new_AGEMA_reg_buffer_10186 ( .C (clk), .D (new_AGEMA_signal_22909), .Q (new_AGEMA_signal_22910) ) ;
    buf_clk new_AGEMA_reg_buffer_10190 ( .C (clk), .D (new_AGEMA_signal_22913), .Q (new_AGEMA_signal_22914) ) ;
    buf_clk new_AGEMA_reg_buffer_10194 ( .C (clk), .D (new_AGEMA_signal_22917), .Q (new_AGEMA_signal_22918) ) ;
    buf_clk new_AGEMA_reg_buffer_10198 ( .C (clk), .D (new_AGEMA_signal_22921), .Q (new_AGEMA_signal_22922) ) ;
    buf_clk new_AGEMA_reg_buffer_10202 ( .C (clk), .D (new_AGEMA_signal_22925), .Q (new_AGEMA_signal_22926) ) ;
    buf_clk new_AGEMA_reg_buffer_10206 ( .C (clk), .D (new_AGEMA_signal_22929), .Q (new_AGEMA_signal_22930) ) ;
    buf_clk new_AGEMA_reg_buffer_10210 ( .C (clk), .D (new_AGEMA_signal_22933), .Q (new_AGEMA_signal_22934) ) ;
    buf_clk new_AGEMA_reg_buffer_10214 ( .C (clk), .D (new_AGEMA_signal_22937), .Q (new_AGEMA_signal_22938) ) ;
    buf_clk new_AGEMA_reg_buffer_10218 ( .C (clk), .D (new_AGEMA_signal_22941), .Q (new_AGEMA_signal_22942) ) ;
    buf_clk new_AGEMA_reg_buffer_10222 ( .C (clk), .D (new_AGEMA_signal_22945), .Q (new_AGEMA_signal_22946) ) ;
    buf_clk new_AGEMA_reg_buffer_10226 ( .C (clk), .D (new_AGEMA_signal_22949), .Q (new_AGEMA_signal_22950) ) ;
    buf_clk new_AGEMA_reg_buffer_10230 ( .C (clk), .D (new_AGEMA_signal_22953), .Q (new_AGEMA_signal_22954) ) ;
    buf_clk new_AGEMA_reg_buffer_10234 ( .C (clk), .D (new_AGEMA_signal_22957), .Q (new_AGEMA_signal_22958) ) ;
    buf_clk new_AGEMA_reg_buffer_10238 ( .C (clk), .D (new_AGEMA_signal_22961), .Q (new_AGEMA_signal_22962) ) ;
    buf_clk new_AGEMA_reg_buffer_10242 ( .C (clk), .D (new_AGEMA_signal_22965), .Q (new_AGEMA_signal_22966) ) ;
    buf_clk new_AGEMA_reg_buffer_10246 ( .C (clk), .D (new_AGEMA_signal_22969), .Q (new_AGEMA_signal_22970) ) ;
    buf_clk new_AGEMA_reg_buffer_10250 ( .C (clk), .D (new_AGEMA_signal_22973), .Q (new_AGEMA_signal_22974) ) ;
    buf_clk new_AGEMA_reg_buffer_10254 ( .C (clk), .D (new_AGEMA_signal_22977), .Q (new_AGEMA_signal_22978) ) ;
    buf_clk new_AGEMA_reg_buffer_10258 ( .C (clk), .D (new_AGEMA_signal_22981), .Q (new_AGEMA_signal_22982) ) ;
    buf_clk new_AGEMA_reg_buffer_10262 ( .C (clk), .D (new_AGEMA_signal_22985), .Q (new_AGEMA_signal_22986) ) ;
    buf_clk new_AGEMA_reg_buffer_10266 ( .C (clk), .D (new_AGEMA_signal_22989), .Q (new_AGEMA_signal_22990) ) ;
    buf_clk new_AGEMA_reg_buffer_10270 ( .C (clk), .D (new_AGEMA_signal_22993), .Q (new_AGEMA_signal_22994) ) ;
    buf_clk new_AGEMA_reg_buffer_10274 ( .C (clk), .D (new_AGEMA_signal_22997), .Q (new_AGEMA_signal_22998) ) ;
    buf_clk new_AGEMA_reg_buffer_10278 ( .C (clk), .D (new_AGEMA_signal_23001), .Q (new_AGEMA_signal_23002) ) ;
    buf_clk new_AGEMA_reg_buffer_10282 ( .C (clk), .D (new_AGEMA_signal_23005), .Q (new_AGEMA_signal_23006) ) ;
    buf_clk new_AGEMA_reg_buffer_10286 ( .C (clk), .D (new_AGEMA_signal_23009), .Q (new_AGEMA_signal_23010) ) ;
    buf_clk new_AGEMA_reg_buffer_10290 ( .C (clk), .D (new_AGEMA_signal_23013), .Q (new_AGEMA_signal_23014) ) ;
    buf_clk new_AGEMA_reg_buffer_10294 ( .C (clk), .D (new_AGEMA_signal_23017), .Q (new_AGEMA_signal_23018) ) ;
    buf_clk new_AGEMA_reg_buffer_10298 ( .C (clk), .D (new_AGEMA_signal_23021), .Q (new_AGEMA_signal_23022) ) ;
    buf_clk new_AGEMA_reg_buffer_10302 ( .C (clk), .D (new_AGEMA_signal_23025), .Q (new_AGEMA_signal_23026) ) ;
    buf_clk new_AGEMA_reg_buffer_10306 ( .C (clk), .D (new_AGEMA_signal_23029), .Q (new_AGEMA_signal_23030) ) ;
    buf_clk new_AGEMA_reg_buffer_10310 ( .C (clk), .D (new_AGEMA_signal_23033), .Q (new_AGEMA_signal_23034) ) ;
    buf_clk new_AGEMA_reg_buffer_10314 ( .C (clk), .D (new_AGEMA_signal_23037), .Q (new_AGEMA_signal_23038) ) ;
    buf_clk new_AGEMA_reg_buffer_10318 ( .C (clk), .D (new_AGEMA_signal_23041), .Q (new_AGEMA_signal_23042) ) ;
    buf_clk new_AGEMA_reg_buffer_10322 ( .C (clk), .D (new_AGEMA_signal_23045), .Q (new_AGEMA_signal_23046) ) ;
    buf_clk new_AGEMA_reg_buffer_10326 ( .C (clk), .D (new_AGEMA_signal_23049), .Q (new_AGEMA_signal_23050) ) ;
    buf_clk new_AGEMA_reg_buffer_10330 ( .C (clk), .D (new_AGEMA_signal_23053), .Q (new_AGEMA_signal_23054) ) ;
    buf_clk new_AGEMA_reg_buffer_10334 ( .C (clk), .D (new_AGEMA_signal_23057), .Q (new_AGEMA_signal_23058) ) ;
    buf_clk new_AGEMA_reg_buffer_10338 ( .C (clk), .D (new_AGEMA_signal_23061), .Q (new_AGEMA_signal_23062) ) ;
    buf_clk new_AGEMA_reg_buffer_10342 ( .C (clk), .D (new_AGEMA_signal_23065), .Q (new_AGEMA_signal_23066) ) ;
    buf_clk new_AGEMA_reg_buffer_10346 ( .C (clk), .D (new_AGEMA_signal_23069), .Q (new_AGEMA_signal_23070) ) ;
    buf_clk new_AGEMA_reg_buffer_10350 ( .C (clk), .D (new_AGEMA_signal_23073), .Q (new_AGEMA_signal_23074) ) ;
    buf_clk new_AGEMA_reg_buffer_10354 ( .C (clk), .D (new_AGEMA_signal_23077), .Q (new_AGEMA_signal_23078) ) ;
    buf_clk new_AGEMA_reg_buffer_10358 ( .C (clk), .D (new_AGEMA_signal_23081), .Q (new_AGEMA_signal_23082) ) ;
    buf_clk new_AGEMA_reg_buffer_10362 ( .C (clk), .D (new_AGEMA_signal_23085), .Q (new_AGEMA_signal_23086) ) ;
    buf_clk new_AGEMA_reg_buffer_10366 ( .C (clk), .D (new_AGEMA_signal_23089), .Q (new_AGEMA_signal_23090) ) ;
    buf_clk new_AGEMA_reg_buffer_10370 ( .C (clk), .D (new_AGEMA_signal_23093), .Q (new_AGEMA_signal_23094) ) ;
    buf_clk new_AGEMA_reg_buffer_10374 ( .C (clk), .D (new_AGEMA_signal_23097), .Q (new_AGEMA_signal_23098) ) ;
    buf_clk new_AGEMA_reg_buffer_10378 ( .C (clk), .D (new_AGEMA_signal_23101), .Q (new_AGEMA_signal_23102) ) ;
    buf_clk new_AGEMA_reg_buffer_10382 ( .C (clk), .D (new_AGEMA_signal_23105), .Q (new_AGEMA_signal_23106) ) ;
    buf_clk new_AGEMA_reg_buffer_10386 ( .C (clk), .D (new_AGEMA_signal_23109), .Q (new_AGEMA_signal_23110) ) ;
    buf_clk new_AGEMA_reg_buffer_10390 ( .C (clk), .D (new_AGEMA_signal_23113), .Q (new_AGEMA_signal_23114) ) ;
    buf_clk new_AGEMA_reg_buffer_10394 ( .C (clk), .D (new_AGEMA_signal_23117), .Q (new_AGEMA_signal_23118) ) ;
    buf_clk new_AGEMA_reg_buffer_10398 ( .C (clk), .D (new_AGEMA_signal_23121), .Q (new_AGEMA_signal_23122) ) ;
    buf_clk new_AGEMA_reg_buffer_10402 ( .C (clk), .D (new_AGEMA_signal_23125), .Q (new_AGEMA_signal_23126) ) ;
    buf_clk new_AGEMA_reg_buffer_10406 ( .C (clk), .D (new_AGEMA_signal_23129), .Q (new_AGEMA_signal_23130) ) ;
    buf_clk new_AGEMA_reg_buffer_10410 ( .C (clk), .D (new_AGEMA_signal_23133), .Q (new_AGEMA_signal_23134) ) ;
    buf_clk new_AGEMA_reg_buffer_10414 ( .C (clk), .D (new_AGEMA_signal_23137), .Q (new_AGEMA_signal_23138) ) ;
    buf_clk new_AGEMA_reg_buffer_10418 ( .C (clk), .D (new_AGEMA_signal_23141), .Q (new_AGEMA_signal_23142) ) ;
    buf_clk new_AGEMA_reg_buffer_10422 ( .C (clk), .D (new_AGEMA_signal_23145), .Q (new_AGEMA_signal_23146) ) ;
    buf_clk new_AGEMA_reg_buffer_10426 ( .C (clk), .D (new_AGEMA_signal_23149), .Q (new_AGEMA_signal_23150) ) ;
    buf_clk new_AGEMA_reg_buffer_10430 ( .C (clk), .D (new_AGEMA_signal_23153), .Q (new_AGEMA_signal_23154) ) ;
    buf_clk new_AGEMA_reg_buffer_10434 ( .C (clk), .D (new_AGEMA_signal_23157), .Q (new_AGEMA_signal_23158) ) ;
    buf_clk new_AGEMA_reg_buffer_10438 ( .C (clk), .D (new_AGEMA_signal_23161), .Q (new_AGEMA_signal_23162) ) ;
    buf_clk new_AGEMA_reg_buffer_10442 ( .C (clk), .D (new_AGEMA_signal_23165), .Q (new_AGEMA_signal_23166) ) ;
    buf_clk new_AGEMA_reg_buffer_10446 ( .C (clk), .D (new_AGEMA_signal_23169), .Q (new_AGEMA_signal_23170) ) ;
    buf_clk new_AGEMA_reg_buffer_10450 ( .C (clk), .D (new_AGEMA_signal_23173), .Q (new_AGEMA_signal_23174) ) ;
    buf_clk new_AGEMA_reg_buffer_10454 ( .C (clk), .D (new_AGEMA_signal_23177), .Q (new_AGEMA_signal_23178) ) ;
    buf_clk new_AGEMA_reg_buffer_10458 ( .C (clk), .D (new_AGEMA_signal_23181), .Q (new_AGEMA_signal_23182) ) ;
    buf_clk new_AGEMA_reg_buffer_10462 ( .C (clk), .D (new_AGEMA_signal_23185), .Q (new_AGEMA_signal_23186) ) ;
    buf_clk new_AGEMA_reg_buffer_10466 ( .C (clk), .D (new_AGEMA_signal_23189), .Q (new_AGEMA_signal_23190) ) ;
    buf_clk new_AGEMA_reg_buffer_10470 ( .C (clk), .D (new_AGEMA_signal_23193), .Q (new_AGEMA_signal_23194) ) ;
    buf_clk new_AGEMA_reg_buffer_10474 ( .C (clk), .D (new_AGEMA_signal_23197), .Q (new_AGEMA_signal_23198) ) ;
    buf_clk new_AGEMA_reg_buffer_10478 ( .C (clk), .D (new_AGEMA_signal_23201), .Q (new_AGEMA_signal_23202) ) ;
    buf_clk new_AGEMA_reg_buffer_10482 ( .C (clk), .D (new_AGEMA_signal_23205), .Q (new_AGEMA_signal_23206) ) ;
    buf_clk new_AGEMA_reg_buffer_10486 ( .C (clk), .D (new_AGEMA_signal_23209), .Q (new_AGEMA_signal_23210) ) ;
    buf_clk new_AGEMA_reg_buffer_10490 ( .C (clk), .D (new_AGEMA_signal_23213), .Q (new_AGEMA_signal_23214) ) ;
    buf_clk new_AGEMA_reg_buffer_10494 ( .C (clk), .D (new_AGEMA_signal_23217), .Q (new_AGEMA_signal_23218) ) ;
    buf_clk new_AGEMA_reg_buffer_10498 ( .C (clk), .D (new_AGEMA_signal_23221), .Q (new_AGEMA_signal_23222) ) ;
    buf_clk new_AGEMA_reg_buffer_10502 ( .C (clk), .D (new_AGEMA_signal_23225), .Q (new_AGEMA_signal_23226) ) ;
    buf_clk new_AGEMA_reg_buffer_10506 ( .C (clk), .D (new_AGEMA_signal_23229), .Q (new_AGEMA_signal_23230) ) ;
    buf_clk new_AGEMA_reg_buffer_10510 ( .C (clk), .D (new_AGEMA_signal_23233), .Q (new_AGEMA_signal_23234) ) ;
    buf_clk new_AGEMA_reg_buffer_10514 ( .C (clk), .D (new_AGEMA_signal_23237), .Q (new_AGEMA_signal_23238) ) ;
    buf_clk new_AGEMA_reg_buffer_10518 ( .C (clk), .D (new_AGEMA_signal_23241), .Q (new_AGEMA_signal_23242) ) ;
    buf_clk new_AGEMA_reg_buffer_10522 ( .C (clk), .D (new_AGEMA_signal_23245), .Q (new_AGEMA_signal_23246) ) ;
    buf_clk new_AGEMA_reg_buffer_10526 ( .C (clk), .D (new_AGEMA_signal_23249), .Q (new_AGEMA_signal_23250) ) ;
    buf_clk new_AGEMA_reg_buffer_10530 ( .C (clk), .D (new_AGEMA_signal_23253), .Q (new_AGEMA_signal_23254) ) ;
    buf_clk new_AGEMA_reg_buffer_10534 ( .C (clk), .D (new_AGEMA_signal_23257), .Q (new_AGEMA_signal_23258) ) ;
    buf_clk new_AGEMA_reg_buffer_10538 ( .C (clk), .D (new_AGEMA_signal_23261), .Q (new_AGEMA_signal_23262) ) ;
    buf_clk new_AGEMA_reg_buffer_10542 ( .C (clk), .D (new_AGEMA_signal_23265), .Q (new_AGEMA_signal_23266) ) ;
    buf_clk new_AGEMA_reg_buffer_10546 ( .C (clk), .D (new_AGEMA_signal_23269), .Q (new_AGEMA_signal_23270) ) ;
    buf_clk new_AGEMA_reg_buffer_10550 ( .C (clk), .D (new_AGEMA_signal_23273), .Q (new_AGEMA_signal_23274) ) ;
    buf_clk new_AGEMA_reg_buffer_10554 ( .C (clk), .D (new_AGEMA_signal_23277), .Q (new_AGEMA_signal_23278) ) ;
    buf_clk new_AGEMA_reg_buffer_10558 ( .C (clk), .D (new_AGEMA_signal_23281), .Q (new_AGEMA_signal_23282) ) ;
    buf_clk new_AGEMA_reg_buffer_10562 ( .C (clk), .D (new_AGEMA_signal_23285), .Q (new_AGEMA_signal_23286) ) ;
    buf_clk new_AGEMA_reg_buffer_10566 ( .C (clk), .D (new_AGEMA_signal_23289), .Q (new_AGEMA_signal_23290) ) ;
    buf_clk new_AGEMA_reg_buffer_10570 ( .C (clk), .D (new_AGEMA_signal_23293), .Q (new_AGEMA_signal_23294) ) ;
    buf_clk new_AGEMA_reg_buffer_10574 ( .C (clk), .D (new_AGEMA_signal_23297), .Q (new_AGEMA_signal_23298) ) ;
    buf_clk new_AGEMA_reg_buffer_10578 ( .C (clk), .D (new_AGEMA_signal_23301), .Q (new_AGEMA_signal_23302) ) ;
    buf_clk new_AGEMA_reg_buffer_10582 ( .C (clk), .D (new_AGEMA_signal_23305), .Q (new_AGEMA_signal_23306) ) ;
    buf_clk new_AGEMA_reg_buffer_10586 ( .C (clk), .D (new_AGEMA_signal_23309), .Q (new_AGEMA_signal_23310) ) ;
    buf_clk new_AGEMA_reg_buffer_10590 ( .C (clk), .D (new_AGEMA_signal_23313), .Q (new_AGEMA_signal_23314) ) ;
    buf_clk new_AGEMA_reg_buffer_10594 ( .C (clk), .D (new_AGEMA_signal_23317), .Q (new_AGEMA_signal_23318) ) ;
    buf_clk new_AGEMA_reg_buffer_10598 ( .C (clk), .D (new_AGEMA_signal_23321), .Q (new_AGEMA_signal_23322) ) ;
    buf_clk new_AGEMA_reg_buffer_10602 ( .C (clk), .D (new_AGEMA_signal_23325), .Q (new_AGEMA_signal_23326) ) ;
    buf_clk new_AGEMA_reg_buffer_10606 ( .C (clk), .D (new_AGEMA_signal_23329), .Q (new_AGEMA_signal_23330) ) ;
    buf_clk new_AGEMA_reg_buffer_10610 ( .C (clk), .D (new_AGEMA_signal_23333), .Q (new_AGEMA_signal_23334) ) ;
    buf_clk new_AGEMA_reg_buffer_10614 ( .C (clk), .D (new_AGEMA_signal_23337), .Q (new_AGEMA_signal_23338) ) ;
    buf_clk new_AGEMA_reg_buffer_10618 ( .C (clk), .D (new_AGEMA_signal_23341), .Q (new_AGEMA_signal_23342) ) ;
    buf_clk new_AGEMA_reg_buffer_10622 ( .C (clk), .D (new_AGEMA_signal_23345), .Q (new_AGEMA_signal_23346) ) ;
    buf_clk new_AGEMA_reg_buffer_10626 ( .C (clk), .D (new_AGEMA_signal_23349), .Q (new_AGEMA_signal_23350) ) ;
    buf_clk new_AGEMA_reg_buffer_10630 ( .C (clk), .D (new_AGEMA_signal_23353), .Q (new_AGEMA_signal_23354) ) ;
    buf_clk new_AGEMA_reg_buffer_10634 ( .C (clk), .D (new_AGEMA_signal_23357), .Q (new_AGEMA_signal_23358) ) ;
    buf_clk new_AGEMA_reg_buffer_10638 ( .C (clk), .D (new_AGEMA_signal_23361), .Q (new_AGEMA_signal_23362) ) ;
    buf_clk new_AGEMA_reg_buffer_10642 ( .C (clk), .D (new_AGEMA_signal_23365), .Q (new_AGEMA_signal_23366) ) ;
    buf_clk new_AGEMA_reg_buffer_10646 ( .C (clk), .D (new_AGEMA_signal_23369), .Q (new_AGEMA_signal_23370) ) ;
    buf_clk new_AGEMA_reg_buffer_10650 ( .C (clk), .D (new_AGEMA_signal_23373), .Q (new_AGEMA_signal_23374) ) ;
    buf_clk new_AGEMA_reg_buffer_10654 ( .C (clk), .D (new_AGEMA_signal_23377), .Q (new_AGEMA_signal_23378) ) ;
    buf_clk new_AGEMA_reg_buffer_10658 ( .C (clk), .D (new_AGEMA_signal_23381), .Q (new_AGEMA_signal_23382) ) ;
    buf_clk new_AGEMA_reg_buffer_10662 ( .C (clk), .D (new_AGEMA_signal_23385), .Q (new_AGEMA_signal_23386) ) ;
    buf_clk new_AGEMA_reg_buffer_10666 ( .C (clk), .D (new_AGEMA_signal_23389), .Q (new_AGEMA_signal_23390) ) ;
    buf_clk new_AGEMA_reg_buffer_10670 ( .C (clk), .D (new_AGEMA_signal_23393), .Q (new_AGEMA_signal_23394) ) ;
    buf_clk new_AGEMA_reg_buffer_10674 ( .C (clk), .D (new_AGEMA_signal_23397), .Q (new_AGEMA_signal_23398) ) ;
    buf_clk new_AGEMA_reg_buffer_10678 ( .C (clk), .D (new_AGEMA_signal_23401), .Q (new_AGEMA_signal_23402) ) ;
    buf_clk new_AGEMA_reg_buffer_10682 ( .C (clk), .D (new_AGEMA_signal_23405), .Q (new_AGEMA_signal_23406) ) ;
    buf_clk new_AGEMA_reg_buffer_10686 ( .C (clk), .D (new_AGEMA_signal_23409), .Q (new_AGEMA_signal_23410) ) ;
    buf_clk new_AGEMA_reg_buffer_10690 ( .C (clk), .D (new_AGEMA_signal_23413), .Q (new_AGEMA_signal_23414) ) ;
    buf_clk new_AGEMA_reg_buffer_10694 ( .C (clk), .D (new_AGEMA_signal_23417), .Q (new_AGEMA_signal_23418) ) ;
    buf_clk new_AGEMA_reg_buffer_10698 ( .C (clk), .D (new_AGEMA_signal_23421), .Q (new_AGEMA_signal_23422) ) ;
    buf_clk new_AGEMA_reg_buffer_10702 ( .C (clk), .D (new_AGEMA_signal_23425), .Q (new_AGEMA_signal_23426) ) ;
    buf_clk new_AGEMA_reg_buffer_10706 ( .C (clk), .D (new_AGEMA_signal_23429), .Q (new_AGEMA_signal_23430) ) ;
    buf_clk new_AGEMA_reg_buffer_10710 ( .C (clk), .D (new_AGEMA_signal_23433), .Q (new_AGEMA_signal_23434) ) ;
    buf_clk new_AGEMA_reg_buffer_10714 ( .C (clk), .D (new_AGEMA_signal_23437), .Q (new_AGEMA_signal_23438) ) ;
    buf_clk new_AGEMA_reg_buffer_10718 ( .C (clk), .D (new_AGEMA_signal_23441), .Q (new_AGEMA_signal_23442) ) ;
    buf_clk new_AGEMA_reg_buffer_10722 ( .C (clk), .D (new_AGEMA_signal_23445), .Q (new_AGEMA_signal_23446) ) ;
    buf_clk new_AGEMA_reg_buffer_10726 ( .C (clk), .D (new_AGEMA_signal_23449), .Q (new_AGEMA_signal_23450) ) ;
    buf_clk new_AGEMA_reg_buffer_10730 ( .C (clk), .D (new_AGEMA_signal_23453), .Q (new_AGEMA_signal_23454) ) ;
    buf_clk new_AGEMA_reg_buffer_10734 ( .C (clk), .D (new_AGEMA_signal_23457), .Q (new_AGEMA_signal_23458) ) ;
    buf_clk new_AGEMA_reg_buffer_10738 ( .C (clk), .D (new_AGEMA_signal_23461), .Q (new_AGEMA_signal_23462) ) ;
    buf_clk new_AGEMA_reg_buffer_10742 ( .C (clk), .D (new_AGEMA_signal_23465), .Q (new_AGEMA_signal_23466) ) ;
    buf_clk new_AGEMA_reg_buffer_10746 ( .C (clk), .D (new_AGEMA_signal_23469), .Q (new_AGEMA_signal_23470) ) ;
    buf_clk new_AGEMA_reg_buffer_10750 ( .C (clk), .D (new_AGEMA_signal_23473), .Q (new_AGEMA_signal_23474) ) ;
    buf_clk new_AGEMA_reg_buffer_10754 ( .C (clk), .D (new_AGEMA_signal_23477), .Q (new_AGEMA_signal_23478) ) ;
    buf_clk new_AGEMA_reg_buffer_10758 ( .C (clk), .D (new_AGEMA_signal_23481), .Q (new_AGEMA_signal_23482) ) ;
    buf_clk new_AGEMA_reg_buffer_10762 ( .C (clk), .D (new_AGEMA_signal_23485), .Q (new_AGEMA_signal_23486) ) ;
    buf_clk new_AGEMA_reg_buffer_10766 ( .C (clk), .D (new_AGEMA_signal_23489), .Q (new_AGEMA_signal_23490) ) ;
    buf_clk new_AGEMA_reg_buffer_10770 ( .C (clk), .D (new_AGEMA_signal_23493), .Q (new_AGEMA_signal_23494) ) ;
    buf_clk new_AGEMA_reg_buffer_10774 ( .C (clk), .D (new_AGEMA_signal_23497), .Q (new_AGEMA_signal_23498) ) ;
    buf_clk new_AGEMA_reg_buffer_10778 ( .C (clk), .D (new_AGEMA_signal_23501), .Q (new_AGEMA_signal_23502) ) ;
    buf_clk new_AGEMA_reg_buffer_10782 ( .C (clk), .D (new_AGEMA_signal_23505), .Q (new_AGEMA_signal_23506) ) ;
    buf_clk new_AGEMA_reg_buffer_10786 ( .C (clk), .D (new_AGEMA_signal_23509), .Q (new_AGEMA_signal_23510) ) ;
    buf_clk new_AGEMA_reg_buffer_10790 ( .C (clk), .D (new_AGEMA_signal_23513), .Q (new_AGEMA_signal_23514) ) ;
    buf_clk new_AGEMA_reg_buffer_10794 ( .C (clk), .D (new_AGEMA_signal_23517), .Q (new_AGEMA_signal_23518) ) ;
    buf_clk new_AGEMA_reg_buffer_10798 ( .C (clk), .D (new_AGEMA_signal_23521), .Q (new_AGEMA_signal_23522) ) ;
    buf_clk new_AGEMA_reg_buffer_10802 ( .C (clk), .D (new_AGEMA_signal_23525), .Q (new_AGEMA_signal_23526) ) ;
    buf_clk new_AGEMA_reg_buffer_10806 ( .C (clk), .D (new_AGEMA_signal_23529), .Q (new_AGEMA_signal_23530) ) ;
    buf_clk new_AGEMA_reg_buffer_10810 ( .C (clk), .D (new_AGEMA_signal_23533), .Q (new_AGEMA_signal_23534) ) ;
    buf_clk new_AGEMA_reg_buffer_10814 ( .C (clk), .D (new_AGEMA_signal_23537), .Q (new_AGEMA_signal_23538) ) ;
    buf_clk new_AGEMA_reg_buffer_10818 ( .C (clk), .D (new_AGEMA_signal_23541), .Q (new_AGEMA_signal_23542) ) ;
    buf_clk new_AGEMA_reg_buffer_10822 ( .C (clk), .D (new_AGEMA_signal_23545), .Q (new_AGEMA_signal_23546) ) ;
    buf_clk new_AGEMA_reg_buffer_10826 ( .C (clk), .D (new_AGEMA_signal_23549), .Q (new_AGEMA_signal_23550) ) ;
    buf_clk new_AGEMA_reg_buffer_10830 ( .C (clk), .D (new_AGEMA_signal_23553), .Q (new_AGEMA_signal_23554) ) ;
    buf_clk new_AGEMA_reg_buffer_10834 ( .C (clk), .D (new_AGEMA_signal_23557), .Q (new_AGEMA_signal_23558) ) ;
    buf_clk new_AGEMA_reg_buffer_10838 ( .C (clk), .D (new_AGEMA_signal_23561), .Q (new_AGEMA_signal_23562) ) ;
    buf_clk new_AGEMA_reg_buffer_10842 ( .C (clk), .D (new_AGEMA_signal_23565), .Q (new_AGEMA_signal_23566) ) ;
    buf_clk new_AGEMA_reg_buffer_10846 ( .C (clk), .D (new_AGEMA_signal_23569), .Q (new_AGEMA_signal_23570) ) ;
    buf_clk new_AGEMA_reg_buffer_10850 ( .C (clk), .D (new_AGEMA_signal_23573), .Q (new_AGEMA_signal_23574) ) ;
    buf_clk new_AGEMA_reg_buffer_10854 ( .C (clk), .D (new_AGEMA_signal_23577), .Q (new_AGEMA_signal_23578) ) ;
    buf_clk new_AGEMA_reg_buffer_10858 ( .C (clk), .D (new_AGEMA_signal_23581), .Q (new_AGEMA_signal_23582) ) ;
    buf_clk new_AGEMA_reg_buffer_10862 ( .C (clk), .D (new_AGEMA_signal_23585), .Q (new_AGEMA_signal_23586) ) ;
    buf_clk new_AGEMA_reg_buffer_10866 ( .C (clk), .D (new_AGEMA_signal_23589), .Q (new_AGEMA_signal_23590) ) ;
    buf_clk new_AGEMA_reg_buffer_10870 ( .C (clk), .D (new_AGEMA_signal_23593), .Q (new_AGEMA_signal_23594) ) ;
    buf_clk new_AGEMA_reg_buffer_10874 ( .C (clk), .D (new_AGEMA_signal_23597), .Q (new_AGEMA_signal_23598) ) ;
    buf_clk new_AGEMA_reg_buffer_10878 ( .C (clk), .D (new_AGEMA_signal_23601), .Q (new_AGEMA_signal_23602) ) ;
    buf_clk new_AGEMA_reg_buffer_10882 ( .C (clk), .D (new_AGEMA_signal_23605), .Q (new_AGEMA_signal_23606) ) ;
    buf_clk new_AGEMA_reg_buffer_10886 ( .C (clk), .D (new_AGEMA_signal_23609), .Q (new_AGEMA_signal_23610) ) ;
    buf_clk new_AGEMA_reg_buffer_10890 ( .C (clk), .D (new_AGEMA_signal_23613), .Q (new_AGEMA_signal_23614) ) ;
    buf_clk new_AGEMA_reg_buffer_10894 ( .C (clk), .D (new_AGEMA_signal_23617), .Q (new_AGEMA_signal_23618) ) ;
    buf_clk new_AGEMA_reg_buffer_10898 ( .C (clk), .D (new_AGEMA_signal_23621), .Q (new_AGEMA_signal_23622) ) ;
    buf_clk new_AGEMA_reg_buffer_10902 ( .C (clk), .D (new_AGEMA_signal_23625), .Q (new_AGEMA_signal_23626) ) ;
    buf_clk new_AGEMA_reg_buffer_10906 ( .C (clk), .D (new_AGEMA_signal_23629), .Q (new_AGEMA_signal_23630) ) ;
    buf_clk new_AGEMA_reg_buffer_10910 ( .C (clk), .D (new_AGEMA_signal_23633), .Q (new_AGEMA_signal_23634) ) ;
    buf_clk new_AGEMA_reg_buffer_10914 ( .C (clk), .D (new_AGEMA_signal_23637), .Q (new_AGEMA_signal_23638) ) ;
    buf_clk new_AGEMA_reg_buffer_10918 ( .C (clk), .D (new_AGEMA_signal_23641), .Q (new_AGEMA_signal_23642) ) ;
    buf_clk new_AGEMA_reg_buffer_10922 ( .C (clk), .D (new_AGEMA_signal_23645), .Q (new_AGEMA_signal_23646) ) ;
    buf_clk new_AGEMA_reg_buffer_10926 ( .C (clk), .D (new_AGEMA_signal_23649), .Q (new_AGEMA_signal_23650) ) ;
    buf_clk new_AGEMA_reg_buffer_10930 ( .C (clk), .D (new_AGEMA_signal_23653), .Q (new_AGEMA_signal_23654) ) ;
    buf_clk new_AGEMA_reg_buffer_10934 ( .C (clk), .D (new_AGEMA_signal_23657), .Q (new_AGEMA_signal_23658) ) ;
    buf_clk new_AGEMA_reg_buffer_10938 ( .C (clk), .D (new_AGEMA_signal_23661), .Q (new_AGEMA_signal_23662) ) ;
    buf_clk new_AGEMA_reg_buffer_10942 ( .C (clk), .D (new_AGEMA_signal_23665), .Q (new_AGEMA_signal_23666) ) ;
    buf_clk new_AGEMA_reg_buffer_10946 ( .C (clk), .D (new_AGEMA_signal_23669), .Q (new_AGEMA_signal_23670) ) ;
    buf_clk new_AGEMA_reg_buffer_10950 ( .C (clk), .D (new_AGEMA_signal_23673), .Q (new_AGEMA_signal_23674) ) ;
    buf_clk new_AGEMA_reg_buffer_10954 ( .C (clk), .D (new_AGEMA_signal_23677), .Q (new_AGEMA_signal_23678) ) ;
    buf_clk new_AGEMA_reg_buffer_10958 ( .C (clk), .D (new_AGEMA_signal_23681), .Q (new_AGEMA_signal_23682) ) ;
    buf_clk new_AGEMA_reg_buffer_10962 ( .C (clk), .D (new_AGEMA_signal_23685), .Q (new_AGEMA_signal_23686) ) ;
    buf_clk new_AGEMA_reg_buffer_10966 ( .C (clk), .D (new_AGEMA_signal_23689), .Q (new_AGEMA_signal_23690) ) ;
    buf_clk new_AGEMA_reg_buffer_10970 ( .C (clk), .D (new_AGEMA_signal_23693), .Q (new_AGEMA_signal_23694) ) ;
    buf_clk new_AGEMA_reg_buffer_10974 ( .C (clk), .D (new_AGEMA_signal_23697), .Q (new_AGEMA_signal_23698) ) ;
    buf_clk new_AGEMA_reg_buffer_10978 ( .C (clk), .D (new_AGEMA_signal_23701), .Q (new_AGEMA_signal_23702) ) ;
    buf_clk new_AGEMA_reg_buffer_10982 ( .C (clk), .D (new_AGEMA_signal_23705), .Q (new_AGEMA_signal_23706) ) ;
    buf_clk new_AGEMA_reg_buffer_10986 ( .C (clk), .D (new_AGEMA_signal_23709), .Q (new_AGEMA_signal_23710) ) ;
    buf_clk new_AGEMA_reg_buffer_10990 ( .C (clk), .D (new_AGEMA_signal_23713), .Q (new_AGEMA_signal_23714) ) ;
    buf_clk new_AGEMA_reg_buffer_10994 ( .C (clk), .D (new_AGEMA_signal_23717), .Q (new_AGEMA_signal_23718) ) ;
    buf_clk new_AGEMA_reg_buffer_10998 ( .C (clk), .D (new_AGEMA_signal_23721), .Q (new_AGEMA_signal_23722) ) ;
    buf_clk new_AGEMA_reg_buffer_11002 ( .C (clk), .D (new_AGEMA_signal_23725), .Q (new_AGEMA_signal_23726) ) ;
    buf_clk new_AGEMA_reg_buffer_11006 ( .C (clk), .D (new_AGEMA_signal_23729), .Q (new_AGEMA_signal_23730) ) ;
    buf_clk new_AGEMA_reg_buffer_11010 ( .C (clk), .D (new_AGEMA_signal_23733), .Q (new_AGEMA_signal_23734) ) ;
    buf_clk new_AGEMA_reg_buffer_11014 ( .C (clk), .D (new_AGEMA_signal_23737), .Q (new_AGEMA_signal_23738) ) ;
    buf_clk new_AGEMA_reg_buffer_11018 ( .C (clk), .D (new_AGEMA_signal_23741), .Q (new_AGEMA_signal_23742) ) ;
    buf_clk new_AGEMA_reg_buffer_11022 ( .C (clk), .D (new_AGEMA_signal_23745), .Q (new_AGEMA_signal_23746) ) ;
    buf_clk new_AGEMA_reg_buffer_11026 ( .C (clk), .D (new_AGEMA_signal_23749), .Q (new_AGEMA_signal_23750) ) ;
    buf_clk new_AGEMA_reg_buffer_11030 ( .C (clk), .D (new_AGEMA_signal_23753), .Q (new_AGEMA_signal_23754) ) ;
    buf_clk new_AGEMA_reg_buffer_11034 ( .C (clk), .D (new_AGEMA_signal_23757), .Q (new_AGEMA_signal_23758) ) ;
    buf_clk new_AGEMA_reg_buffer_11038 ( .C (clk), .D (new_AGEMA_signal_23761), .Q (new_AGEMA_signal_23762) ) ;
    buf_clk new_AGEMA_reg_buffer_11042 ( .C (clk), .D (new_AGEMA_signal_23765), .Q (new_AGEMA_signal_23766) ) ;
    buf_clk new_AGEMA_reg_buffer_11046 ( .C (clk), .D (new_AGEMA_signal_23769), .Q (new_AGEMA_signal_23770) ) ;
    buf_clk new_AGEMA_reg_buffer_11050 ( .C (clk), .D (new_AGEMA_signal_23773), .Q (new_AGEMA_signal_23774) ) ;
    buf_clk new_AGEMA_reg_buffer_11054 ( .C (clk), .D (new_AGEMA_signal_23777), .Q (new_AGEMA_signal_23778) ) ;
    buf_clk new_AGEMA_reg_buffer_11058 ( .C (clk), .D (new_AGEMA_signal_23781), .Q (new_AGEMA_signal_23782) ) ;
    buf_clk new_AGEMA_reg_buffer_11062 ( .C (clk), .D (new_AGEMA_signal_23785), .Q (new_AGEMA_signal_23786) ) ;
    buf_clk new_AGEMA_reg_buffer_11066 ( .C (clk), .D (new_AGEMA_signal_23789), .Q (new_AGEMA_signal_23790) ) ;
    buf_clk new_AGEMA_reg_buffer_11070 ( .C (clk), .D (new_AGEMA_signal_23793), .Q (new_AGEMA_signal_23794) ) ;
    buf_clk new_AGEMA_reg_buffer_11074 ( .C (clk), .D (new_AGEMA_signal_23797), .Q (new_AGEMA_signal_23798) ) ;
    buf_clk new_AGEMA_reg_buffer_11078 ( .C (clk), .D (new_AGEMA_signal_23801), .Q (new_AGEMA_signal_23802) ) ;
    buf_clk new_AGEMA_reg_buffer_11082 ( .C (clk), .D (new_AGEMA_signal_23805), .Q (new_AGEMA_signal_23806) ) ;
    buf_clk new_AGEMA_reg_buffer_11086 ( .C (clk), .D (new_AGEMA_signal_23809), .Q (new_AGEMA_signal_23810) ) ;
    buf_clk new_AGEMA_reg_buffer_11090 ( .C (clk), .D (new_AGEMA_signal_23813), .Q (new_AGEMA_signal_23814) ) ;
    buf_clk new_AGEMA_reg_buffer_11094 ( .C (clk), .D (new_AGEMA_signal_23817), .Q (new_AGEMA_signal_23818) ) ;
    buf_clk new_AGEMA_reg_buffer_11098 ( .C (clk), .D (new_AGEMA_signal_23821), .Q (new_AGEMA_signal_23822) ) ;
    buf_clk new_AGEMA_reg_buffer_11102 ( .C (clk), .D (new_AGEMA_signal_23825), .Q (new_AGEMA_signal_23826) ) ;
    buf_clk new_AGEMA_reg_buffer_11106 ( .C (clk), .D (new_AGEMA_signal_23829), .Q (new_AGEMA_signal_23830) ) ;
    buf_clk new_AGEMA_reg_buffer_11110 ( .C (clk), .D (new_AGEMA_signal_23833), .Q (new_AGEMA_signal_23834) ) ;
    buf_clk new_AGEMA_reg_buffer_11114 ( .C (clk), .D (new_AGEMA_signal_23837), .Q (new_AGEMA_signal_23838) ) ;
    buf_clk new_AGEMA_reg_buffer_11118 ( .C (clk), .D (new_AGEMA_signal_23841), .Q (new_AGEMA_signal_23842) ) ;
    buf_clk new_AGEMA_reg_buffer_11122 ( .C (clk), .D (new_AGEMA_signal_23845), .Q (new_AGEMA_signal_23846) ) ;
    buf_clk new_AGEMA_reg_buffer_11126 ( .C (clk), .D (new_AGEMA_signal_23849), .Q (new_AGEMA_signal_23850) ) ;
    buf_clk new_AGEMA_reg_buffer_11130 ( .C (clk), .D (new_AGEMA_signal_23853), .Q (new_AGEMA_signal_23854) ) ;
    buf_clk new_AGEMA_reg_buffer_11134 ( .C (clk), .D (new_AGEMA_signal_23857), .Q (new_AGEMA_signal_23858) ) ;
    buf_clk new_AGEMA_reg_buffer_11138 ( .C (clk), .D (new_AGEMA_signal_23861), .Q (new_AGEMA_signal_23862) ) ;
    buf_clk new_AGEMA_reg_buffer_11142 ( .C (clk), .D (new_AGEMA_signal_23865), .Q (new_AGEMA_signal_23866) ) ;
    buf_clk new_AGEMA_reg_buffer_11146 ( .C (clk), .D (new_AGEMA_signal_23869), .Q (new_AGEMA_signal_23870) ) ;
    buf_clk new_AGEMA_reg_buffer_11150 ( .C (clk), .D (new_AGEMA_signal_23873), .Q (new_AGEMA_signal_23874) ) ;
    buf_clk new_AGEMA_reg_buffer_11154 ( .C (clk), .D (new_AGEMA_signal_23877), .Q (new_AGEMA_signal_23878) ) ;
    buf_clk new_AGEMA_reg_buffer_11158 ( .C (clk), .D (new_AGEMA_signal_23881), .Q (new_AGEMA_signal_23882) ) ;
    buf_clk new_AGEMA_reg_buffer_11162 ( .C (clk), .D (new_AGEMA_signal_23885), .Q (new_AGEMA_signal_23886) ) ;
    buf_clk new_AGEMA_reg_buffer_11166 ( .C (clk), .D (new_AGEMA_signal_23889), .Q (new_AGEMA_signal_23890) ) ;
    buf_clk new_AGEMA_reg_buffer_11170 ( .C (clk), .D (new_AGEMA_signal_23893), .Q (new_AGEMA_signal_23894) ) ;
    buf_clk new_AGEMA_reg_buffer_11174 ( .C (clk), .D (new_AGEMA_signal_23897), .Q (new_AGEMA_signal_23898) ) ;
    buf_clk new_AGEMA_reg_buffer_11178 ( .C (clk), .D (new_AGEMA_signal_23901), .Q (new_AGEMA_signal_23902) ) ;
    buf_clk new_AGEMA_reg_buffer_11182 ( .C (clk), .D (new_AGEMA_signal_23905), .Q (new_AGEMA_signal_23906) ) ;
    buf_clk new_AGEMA_reg_buffer_11186 ( .C (clk), .D (new_AGEMA_signal_23909), .Q (new_AGEMA_signal_23910) ) ;
    buf_clk new_AGEMA_reg_buffer_11190 ( .C (clk), .D (new_AGEMA_signal_23913), .Q (new_AGEMA_signal_23914) ) ;
    buf_clk new_AGEMA_reg_buffer_11194 ( .C (clk), .D (new_AGEMA_signal_23917), .Q (new_AGEMA_signal_23918) ) ;
    buf_clk new_AGEMA_reg_buffer_11198 ( .C (clk), .D (new_AGEMA_signal_23921), .Q (new_AGEMA_signal_23922) ) ;
    buf_clk new_AGEMA_reg_buffer_11202 ( .C (clk), .D (new_AGEMA_signal_23925), .Q (new_AGEMA_signal_23926) ) ;
    buf_clk new_AGEMA_reg_buffer_11206 ( .C (clk), .D (new_AGEMA_signal_23929), .Q (new_AGEMA_signal_23930) ) ;
    buf_clk new_AGEMA_reg_buffer_11210 ( .C (clk), .D (new_AGEMA_signal_23933), .Q (new_AGEMA_signal_23934) ) ;
    buf_clk new_AGEMA_reg_buffer_11214 ( .C (clk), .D (new_AGEMA_signal_23937), .Q (new_AGEMA_signal_23938) ) ;
    buf_clk new_AGEMA_reg_buffer_11218 ( .C (clk), .D (new_AGEMA_signal_23941), .Q (new_AGEMA_signal_23942) ) ;
    buf_clk new_AGEMA_reg_buffer_11222 ( .C (clk), .D (new_AGEMA_signal_23945), .Q (new_AGEMA_signal_23946) ) ;
    buf_clk new_AGEMA_reg_buffer_11226 ( .C (clk), .D (new_AGEMA_signal_23949), .Q (new_AGEMA_signal_23950) ) ;
    buf_clk new_AGEMA_reg_buffer_11230 ( .C (clk), .D (new_AGEMA_signal_23953), .Q (new_AGEMA_signal_23954) ) ;
    buf_clk new_AGEMA_reg_buffer_11234 ( .C (clk), .D (new_AGEMA_signal_23957), .Q (new_AGEMA_signal_23958) ) ;
    buf_clk new_AGEMA_reg_buffer_11238 ( .C (clk), .D (new_AGEMA_signal_23961), .Q (new_AGEMA_signal_23962) ) ;
    buf_clk new_AGEMA_reg_buffer_11242 ( .C (clk), .D (new_AGEMA_signal_23965), .Q (new_AGEMA_signal_23966) ) ;
    buf_clk new_AGEMA_reg_buffer_11246 ( .C (clk), .D (new_AGEMA_signal_23969), .Q (new_AGEMA_signal_23970) ) ;
    buf_clk new_AGEMA_reg_buffer_11250 ( .C (clk), .D (new_AGEMA_signal_23973), .Q (new_AGEMA_signal_23974) ) ;
    buf_clk new_AGEMA_reg_buffer_11254 ( .C (clk), .D (new_AGEMA_signal_23977), .Q (new_AGEMA_signal_23978) ) ;
    buf_clk new_AGEMA_reg_buffer_11258 ( .C (clk), .D (new_AGEMA_signal_23981), .Q (new_AGEMA_signal_23982) ) ;
    buf_clk new_AGEMA_reg_buffer_11262 ( .C (clk), .D (new_AGEMA_signal_23985), .Q (new_AGEMA_signal_23986) ) ;
    buf_clk new_AGEMA_reg_buffer_11266 ( .C (clk), .D (new_AGEMA_signal_23989), .Q (new_AGEMA_signal_23990) ) ;
    buf_clk new_AGEMA_reg_buffer_11270 ( .C (clk), .D (new_AGEMA_signal_23993), .Q (new_AGEMA_signal_23994) ) ;
    buf_clk new_AGEMA_reg_buffer_11274 ( .C (clk), .D (new_AGEMA_signal_23997), .Q (new_AGEMA_signal_23998) ) ;
    buf_clk new_AGEMA_reg_buffer_11278 ( .C (clk), .D (new_AGEMA_signal_24001), .Q (new_AGEMA_signal_24002) ) ;
    buf_clk new_AGEMA_reg_buffer_11282 ( .C (clk), .D (new_AGEMA_signal_24005), .Q (new_AGEMA_signal_24006) ) ;
    buf_clk new_AGEMA_reg_buffer_11286 ( .C (clk), .D (new_AGEMA_signal_24009), .Q (new_AGEMA_signal_24010) ) ;
    buf_clk new_AGEMA_reg_buffer_11290 ( .C (clk), .D (new_AGEMA_signal_24013), .Q (new_AGEMA_signal_24014) ) ;
    buf_clk new_AGEMA_reg_buffer_11294 ( .C (clk), .D (new_AGEMA_signal_24017), .Q (new_AGEMA_signal_24018) ) ;
    buf_clk new_AGEMA_reg_buffer_11298 ( .C (clk), .D (new_AGEMA_signal_24021), .Q (new_AGEMA_signal_24022) ) ;
    buf_clk new_AGEMA_reg_buffer_11302 ( .C (clk), .D (new_AGEMA_signal_24025), .Q (new_AGEMA_signal_24026) ) ;
    buf_clk new_AGEMA_reg_buffer_11306 ( .C (clk), .D (new_AGEMA_signal_24029), .Q (new_AGEMA_signal_24030) ) ;
    buf_clk new_AGEMA_reg_buffer_11310 ( .C (clk), .D (new_AGEMA_signal_24033), .Q (new_AGEMA_signal_24034) ) ;
    buf_clk new_AGEMA_reg_buffer_11314 ( .C (clk), .D (new_AGEMA_signal_24037), .Q (new_AGEMA_signal_24038) ) ;
    buf_clk new_AGEMA_reg_buffer_11318 ( .C (clk), .D (new_AGEMA_signal_24041), .Q (new_AGEMA_signal_24042) ) ;
    buf_clk new_AGEMA_reg_buffer_11322 ( .C (clk), .D (new_AGEMA_signal_24045), .Q (new_AGEMA_signal_24046) ) ;
    buf_clk new_AGEMA_reg_buffer_11326 ( .C (clk), .D (new_AGEMA_signal_24049), .Q (new_AGEMA_signal_24050) ) ;
    buf_clk new_AGEMA_reg_buffer_11330 ( .C (clk), .D (new_AGEMA_signal_24053), .Q (new_AGEMA_signal_24054) ) ;
    buf_clk new_AGEMA_reg_buffer_11334 ( .C (clk), .D (new_AGEMA_signal_24057), .Q (new_AGEMA_signal_24058) ) ;
    buf_clk new_AGEMA_reg_buffer_11338 ( .C (clk), .D (new_AGEMA_signal_24061), .Q (new_AGEMA_signal_24062) ) ;
    buf_clk new_AGEMA_reg_buffer_11342 ( .C (clk), .D (new_AGEMA_signal_24065), .Q (new_AGEMA_signal_24066) ) ;
    buf_clk new_AGEMA_reg_buffer_11346 ( .C (clk), .D (new_AGEMA_signal_24069), .Q (new_AGEMA_signal_24070) ) ;
    buf_clk new_AGEMA_reg_buffer_11350 ( .C (clk), .D (new_AGEMA_signal_24073), .Q (new_AGEMA_signal_24074) ) ;
    buf_clk new_AGEMA_reg_buffer_11354 ( .C (clk), .D (new_AGEMA_signal_24077), .Q (new_AGEMA_signal_24078) ) ;
    buf_clk new_AGEMA_reg_buffer_11358 ( .C (clk), .D (new_AGEMA_signal_24081), .Q (new_AGEMA_signal_24082) ) ;
    buf_clk new_AGEMA_reg_buffer_11362 ( .C (clk), .D (new_AGEMA_signal_24085), .Q (new_AGEMA_signal_24086) ) ;
    buf_clk new_AGEMA_reg_buffer_11366 ( .C (clk), .D (new_AGEMA_signal_24089), .Q (new_AGEMA_signal_24090) ) ;
    buf_clk new_AGEMA_reg_buffer_11370 ( .C (clk), .D (new_AGEMA_signal_24093), .Q (new_AGEMA_signal_24094) ) ;
    buf_clk new_AGEMA_reg_buffer_11374 ( .C (clk), .D (new_AGEMA_signal_24097), .Q (new_AGEMA_signal_24098) ) ;
    buf_clk new_AGEMA_reg_buffer_11378 ( .C (clk), .D (new_AGEMA_signal_24101), .Q (new_AGEMA_signal_24102) ) ;
    buf_clk new_AGEMA_reg_buffer_11382 ( .C (clk), .D (new_AGEMA_signal_24105), .Q (new_AGEMA_signal_24106) ) ;
    buf_clk new_AGEMA_reg_buffer_11386 ( .C (clk), .D (new_AGEMA_signal_24109), .Q (new_AGEMA_signal_24110) ) ;
    buf_clk new_AGEMA_reg_buffer_11390 ( .C (clk), .D (new_AGEMA_signal_24113), .Q (new_AGEMA_signal_24114) ) ;
    buf_clk new_AGEMA_reg_buffer_11394 ( .C (clk), .D (new_AGEMA_signal_24117), .Q (new_AGEMA_signal_24118) ) ;
    buf_clk new_AGEMA_reg_buffer_11398 ( .C (clk), .D (new_AGEMA_signal_24121), .Q (new_AGEMA_signal_24122) ) ;
    buf_clk new_AGEMA_reg_buffer_11402 ( .C (clk), .D (new_AGEMA_signal_24125), .Q (new_AGEMA_signal_24126) ) ;
    buf_clk new_AGEMA_reg_buffer_11406 ( .C (clk), .D (new_AGEMA_signal_24129), .Q (new_AGEMA_signal_24130) ) ;
    buf_clk new_AGEMA_reg_buffer_11410 ( .C (clk), .D (new_AGEMA_signal_24133), .Q (new_AGEMA_signal_24134) ) ;
    buf_clk new_AGEMA_reg_buffer_11414 ( .C (clk), .D (new_AGEMA_signal_24137), .Q (new_AGEMA_signal_24138) ) ;
    buf_clk new_AGEMA_reg_buffer_11418 ( .C (clk), .D (new_AGEMA_signal_24141), .Q (new_AGEMA_signal_24142) ) ;
    buf_clk new_AGEMA_reg_buffer_11422 ( .C (clk), .D (new_AGEMA_signal_24145), .Q (new_AGEMA_signal_24146) ) ;
    buf_clk new_AGEMA_reg_buffer_11426 ( .C (clk), .D (new_AGEMA_signal_24149), .Q (new_AGEMA_signal_24150) ) ;
    buf_clk new_AGEMA_reg_buffer_11430 ( .C (clk), .D (new_AGEMA_signal_24153), .Q (new_AGEMA_signal_24154) ) ;
    buf_clk new_AGEMA_reg_buffer_11434 ( .C (clk), .D (new_AGEMA_signal_24157), .Q (new_AGEMA_signal_24158) ) ;
    buf_clk new_AGEMA_reg_buffer_11438 ( .C (clk), .D (new_AGEMA_signal_24161), .Q (new_AGEMA_signal_24162) ) ;
    buf_clk new_AGEMA_reg_buffer_11442 ( .C (clk), .D (new_AGEMA_signal_24165), .Q (new_AGEMA_signal_24166) ) ;
    buf_clk new_AGEMA_reg_buffer_11446 ( .C (clk), .D (new_AGEMA_signal_24169), .Q (new_AGEMA_signal_24170) ) ;
    buf_clk new_AGEMA_reg_buffer_11450 ( .C (clk), .D (new_AGEMA_signal_24173), .Q (new_AGEMA_signal_24174) ) ;
    buf_clk new_AGEMA_reg_buffer_11454 ( .C (clk), .D (new_AGEMA_signal_24177), .Q (new_AGEMA_signal_24178) ) ;
    buf_clk new_AGEMA_reg_buffer_11458 ( .C (clk), .D (new_AGEMA_signal_24181), .Q (new_AGEMA_signal_24182) ) ;
    buf_clk new_AGEMA_reg_buffer_11462 ( .C (clk), .D (new_AGEMA_signal_24185), .Q (new_AGEMA_signal_24186) ) ;
    buf_clk new_AGEMA_reg_buffer_11466 ( .C (clk), .D (new_AGEMA_signal_24189), .Q (new_AGEMA_signal_24190) ) ;
    buf_clk new_AGEMA_reg_buffer_11470 ( .C (clk), .D (new_AGEMA_signal_24193), .Q (new_AGEMA_signal_24194) ) ;
    buf_clk new_AGEMA_reg_buffer_11474 ( .C (clk), .D (new_AGEMA_signal_24197), .Q (new_AGEMA_signal_24198) ) ;
    buf_clk new_AGEMA_reg_buffer_11478 ( .C (clk), .D (new_AGEMA_signal_24201), .Q (new_AGEMA_signal_24202) ) ;
    buf_clk new_AGEMA_reg_buffer_11482 ( .C (clk), .D (new_AGEMA_signal_24205), .Q (new_AGEMA_signal_24206) ) ;
    buf_clk new_AGEMA_reg_buffer_11486 ( .C (clk), .D (new_AGEMA_signal_24209), .Q (new_AGEMA_signal_24210) ) ;
    buf_clk new_AGEMA_reg_buffer_11490 ( .C (clk), .D (new_AGEMA_signal_24213), .Q (new_AGEMA_signal_24214) ) ;
    buf_clk new_AGEMA_reg_buffer_11494 ( .C (clk), .D (new_AGEMA_signal_24217), .Q (new_AGEMA_signal_24218) ) ;
    buf_clk new_AGEMA_reg_buffer_11498 ( .C (clk), .D (new_AGEMA_signal_24221), .Q (new_AGEMA_signal_24222) ) ;
    buf_clk new_AGEMA_reg_buffer_11502 ( .C (clk), .D (new_AGEMA_signal_24225), .Q (new_AGEMA_signal_24226) ) ;
    buf_clk new_AGEMA_reg_buffer_11506 ( .C (clk), .D (new_AGEMA_signal_24229), .Q (new_AGEMA_signal_24230) ) ;
    buf_clk new_AGEMA_reg_buffer_11510 ( .C (clk), .D (new_AGEMA_signal_24233), .Q (new_AGEMA_signal_24234) ) ;
    buf_clk new_AGEMA_reg_buffer_11514 ( .C (clk), .D (new_AGEMA_signal_24237), .Q (new_AGEMA_signal_24238) ) ;
    buf_clk new_AGEMA_reg_buffer_11518 ( .C (clk), .D (new_AGEMA_signal_24241), .Q (new_AGEMA_signal_24242) ) ;
    buf_clk new_AGEMA_reg_buffer_11522 ( .C (clk), .D (new_AGEMA_signal_24245), .Q (new_AGEMA_signal_24246) ) ;
    buf_clk new_AGEMA_reg_buffer_11526 ( .C (clk), .D (new_AGEMA_signal_24249), .Q (new_AGEMA_signal_24250) ) ;
    buf_clk new_AGEMA_reg_buffer_11530 ( .C (clk), .D (new_AGEMA_signal_24253), .Q (new_AGEMA_signal_24254) ) ;
    buf_clk new_AGEMA_reg_buffer_11534 ( .C (clk), .D (new_AGEMA_signal_24257), .Q (new_AGEMA_signal_24258) ) ;
    buf_clk new_AGEMA_reg_buffer_11538 ( .C (clk), .D (new_AGEMA_signal_24261), .Q (new_AGEMA_signal_24262) ) ;
    buf_clk new_AGEMA_reg_buffer_11542 ( .C (clk), .D (new_AGEMA_signal_24265), .Q (new_AGEMA_signal_24266) ) ;
    buf_clk new_AGEMA_reg_buffer_11546 ( .C (clk), .D (new_AGEMA_signal_24269), .Q (new_AGEMA_signal_24270) ) ;
    buf_clk new_AGEMA_reg_buffer_11550 ( .C (clk), .D (new_AGEMA_signal_24273), .Q (new_AGEMA_signal_24274) ) ;
    buf_clk new_AGEMA_reg_buffer_11554 ( .C (clk), .D (new_AGEMA_signal_24277), .Q (new_AGEMA_signal_24278) ) ;
    buf_clk new_AGEMA_reg_buffer_11558 ( .C (clk), .D (new_AGEMA_signal_24281), .Q (new_AGEMA_signal_24282) ) ;
    buf_clk new_AGEMA_reg_buffer_11562 ( .C (clk), .D (new_AGEMA_signal_24285), .Q (new_AGEMA_signal_24286) ) ;
    buf_clk new_AGEMA_reg_buffer_11566 ( .C (clk), .D (new_AGEMA_signal_24289), .Q (new_AGEMA_signal_24290) ) ;
    buf_clk new_AGEMA_reg_buffer_11570 ( .C (clk), .D (new_AGEMA_signal_24293), .Q (new_AGEMA_signal_24294) ) ;
    buf_clk new_AGEMA_reg_buffer_11574 ( .C (clk), .D (new_AGEMA_signal_24297), .Q (new_AGEMA_signal_24298) ) ;
    buf_clk new_AGEMA_reg_buffer_11578 ( .C (clk), .D (new_AGEMA_signal_24301), .Q (new_AGEMA_signal_24302) ) ;
    buf_clk new_AGEMA_reg_buffer_11582 ( .C (clk), .D (new_AGEMA_signal_24305), .Q (new_AGEMA_signal_24306) ) ;
    buf_clk new_AGEMA_reg_buffer_11586 ( .C (clk), .D (new_AGEMA_signal_24309), .Q (new_AGEMA_signal_24310) ) ;
    buf_clk new_AGEMA_reg_buffer_11590 ( .C (clk), .D (new_AGEMA_signal_24313), .Q (new_AGEMA_signal_24314) ) ;
    buf_clk new_AGEMA_reg_buffer_11594 ( .C (clk), .D (new_AGEMA_signal_24317), .Q (new_AGEMA_signal_24318) ) ;
    buf_clk new_AGEMA_reg_buffer_11598 ( .C (clk), .D (new_AGEMA_signal_24321), .Q (new_AGEMA_signal_24322) ) ;
    buf_clk new_AGEMA_reg_buffer_11602 ( .C (clk), .D (new_AGEMA_signal_24325), .Q (new_AGEMA_signal_24326) ) ;
    buf_clk new_AGEMA_reg_buffer_11606 ( .C (clk), .D (new_AGEMA_signal_24329), .Q (new_AGEMA_signal_24330) ) ;
    buf_clk new_AGEMA_reg_buffer_11610 ( .C (clk), .D (new_AGEMA_signal_24333), .Q (new_AGEMA_signal_24334) ) ;
    buf_clk new_AGEMA_reg_buffer_11614 ( .C (clk), .D (new_AGEMA_signal_24337), .Q (new_AGEMA_signal_24338) ) ;
    buf_clk new_AGEMA_reg_buffer_11618 ( .C (clk), .D (new_AGEMA_signal_24341), .Q (new_AGEMA_signal_24342) ) ;
    buf_clk new_AGEMA_reg_buffer_11622 ( .C (clk), .D (new_AGEMA_signal_24345), .Q (new_AGEMA_signal_24346) ) ;
    buf_clk new_AGEMA_reg_buffer_11626 ( .C (clk), .D (new_AGEMA_signal_24349), .Q (new_AGEMA_signal_24350) ) ;
    buf_clk new_AGEMA_reg_buffer_11630 ( .C (clk), .D (new_AGEMA_signal_24353), .Q (new_AGEMA_signal_24354) ) ;
    buf_clk new_AGEMA_reg_buffer_11634 ( .C (clk), .D (new_AGEMA_signal_24357), .Q (new_AGEMA_signal_24358) ) ;
    buf_clk new_AGEMA_reg_buffer_11638 ( .C (clk), .D (new_AGEMA_signal_24361), .Q (new_AGEMA_signal_24362) ) ;
    buf_clk new_AGEMA_reg_buffer_11642 ( .C (clk), .D (new_AGEMA_signal_24365), .Q (new_AGEMA_signal_24366) ) ;
    buf_clk new_AGEMA_reg_buffer_11646 ( .C (clk), .D (new_AGEMA_signal_24369), .Q (new_AGEMA_signal_24370) ) ;
    buf_clk new_AGEMA_reg_buffer_11650 ( .C (clk), .D (new_AGEMA_signal_24373), .Q (new_AGEMA_signal_24374) ) ;
    buf_clk new_AGEMA_reg_buffer_11654 ( .C (clk), .D (new_AGEMA_signal_24377), .Q (new_AGEMA_signal_24378) ) ;
    buf_clk new_AGEMA_reg_buffer_11658 ( .C (clk), .D (new_AGEMA_signal_24381), .Q (new_AGEMA_signal_24382) ) ;
    buf_clk new_AGEMA_reg_buffer_11662 ( .C (clk), .D (new_AGEMA_signal_24385), .Q (new_AGEMA_signal_24386) ) ;
    buf_clk new_AGEMA_reg_buffer_11666 ( .C (clk), .D (new_AGEMA_signal_24389), .Q (new_AGEMA_signal_24390) ) ;
    buf_clk new_AGEMA_reg_buffer_11670 ( .C (clk), .D (new_AGEMA_signal_24393), .Q (new_AGEMA_signal_24394) ) ;
    buf_clk new_AGEMA_reg_buffer_11674 ( .C (clk), .D (new_AGEMA_signal_24397), .Q (new_AGEMA_signal_24398) ) ;
    buf_clk new_AGEMA_reg_buffer_11678 ( .C (clk), .D (new_AGEMA_signal_24401), .Q (new_AGEMA_signal_24402) ) ;
    buf_clk new_AGEMA_reg_buffer_11682 ( .C (clk), .D (new_AGEMA_signal_24405), .Q (new_AGEMA_signal_24406) ) ;
    buf_clk new_AGEMA_reg_buffer_11686 ( .C (clk), .D (new_AGEMA_signal_24409), .Q (new_AGEMA_signal_24410) ) ;
    buf_clk new_AGEMA_reg_buffer_11690 ( .C (clk), .D (new_AGEMA_signal_24413), .Q (new_AGEMA_signal_24414) ) ;
    buf_clk new_AGEMA_reg_buffer_11694 ( .C (clk), .D (new_AGEMA_signal_24417), .Q (new_AGEMA_signal_24418) ) ;
    buf_clk new_AGEMA_reg_buffer_11698 ( .C (clk), .D (new_AGEMA_signal_24421), .Q (new_AGEMA_signal_24422) ) ;
    buf_clk new_AGEMA_reg_buffer_11702 ( .C (clk), .D (new_AGEMA_signal_24425), .Q (new_AGEMA_signal_24426) ) ;
    buf_clk new_AGEMA_reg_buffer_11706 ( .C (clk), .D (new_AGEMA_signal_24429), .Q (new_AGEMA_signal_24430) ) ;
    buf_clk new_AGEMA_reg_buffer_11710 ( .C (clk), .D (new_AGEMA_signal_24433), .Q (new_AGEMA_signal_24434) ) ;
    buf_clk new_AGEMA_reg_buffer_11714 ( .C (clk), .D (new_AGEMA_signal_24437), .Q (new_AGEMA_signal_24438) ) ;
    buf_clk new_AGEMA_reg_buffer_11718 ( .C (clk), .D (new_AGEMA_signal_24441), .Q (new_AGEMA_signal_24442) ) ;
    buf_clk new_AGEMA_reg_buffer_11722 ( .C (clk), .D (new_AGEMA_signal_24445), .Q (new_AGEMA_signal_24446) ) ;
    buf_clk new_AGEMA_reg_buffer_11726 ( .C (clk), .D (new_AGEMA_signal_24449), .Q (new_AGEMA_signal_24450) ) ;
    buf_clk new_AGEMA_reg_buffer_11730 ( .C (clk), .D (new_AGEMA_signal_24453), .Q (new_AGEMA_signal_24454) ) ;
    buf_clk new_AGEMA_reg_buffer_11734 ( .C (clk), .D (new_AGEMA_signal_24457), .Q (new_AGEMA_signal_24458) ) ;
    buf_clk new_AGEMA_reg_buffer_11738 ( .C (clk), .D (new_AGEMA_signal_24461), .Q (new_AGEMA_signal_24462) ) ;
    buf_clk new_AGEMA_reg_buffer_11742 ( .C (clk), .D (new_AGEMA_signal_24465), .Q (new_AGEMA_signal_24466) ) ;
    buf_clk new_AGEMA_reg_buffer_11746 ( .C (clk), .D (new_AGEMA_signal_24469), .Q (new_AGEMA_signal_24470) ) ;
    buf_clk new_AGEMA_reg_buffer_11750 ( .C (clk), .D (new_AGEMA_signal_24473), .Q (new_AGEMA_signal_24474) ) ;
    buf_clk new_AGEMA_reg_buffer_11754 ( .C (clk), .D (new_AGEMA_signal_24477), .Q (new_AGEMA_signal_24478) ) ;
    buf_clk new_AGEMA_reg_buffer_11758 ( .C (clk), .D (new_AGEMA_signal_24481), .Q (new_AGEMA_signal_24482) ) ;
    buf_clk new_AGEMA_reg_buffer_11762 ( .C (clk), .D (new_AGEMA_signal_24485), .Q (new_AGEMA_signal_24486) ) ;
    buf_clk new_AGEMA_reg_buffer_11766 ( .C (clk), .D (new_AGEMA_signal_24489), .Q (new_AGEMA_signal_24490) ) ;
    buf_clk new_AGEMA_reg_buffer_11770 ( .C (clk), .D (new_AGEMA_signal_24493), .Q (new_AGEMA_signal_24494) ) ;
    buf_clk new_AGEMA_reg_buffer_11774 ( .C (clk), .D (new_AGEMA_signal_24497), .Q (new_AGEMA_signal_24498) ) ;
    buf_clk new_AGEMA_reg_buffer_11778 ( .C (clk), .D (new_AGEMA_signal_24501), .Q (new_AGEMA_signal_24502) ) ;
    buf_clk new_AGEMA_reg_buffer_11782 ( .C (clk), .D (new_AGEMA_signal_24505), .Q (new_AGEMA_signal_24506) ) ;
    buf_clk new_AGEMA_reg_buffer_11786 ( .C (clk), .D (new_AGEMA_signal_24509), .Q (new_AGEMA_signal_24510) ) ;
    buf_clk new_AGEMA_reg_buffer_11790 ( .C (clk), .D (new_AGEMA_signal_24513), .Q (new_AGEMA_signal_24514) ) ;
    buf_clk new_AGEMA_reg_buffer_11794 ( .C (clk), .D (new_AGEMA_signal_24517), .Q (new_AGEMA_signal_24518) ) ;
    buf_clk new_AGEMA_reg_buffer_11798 ( .C (clk), .D (new_AGEMA_signal_24521), .Q (new_AGEMA_signal_24522) ) ;
    buf_clk new_AGEMA_reg_buffer_11802 ( .C (clk), .D (new_AGEMA_signal_24525), .Q (new_AGEMA_signal_24526) ) ;
    buf_clk new_AGEMA_reg_buffer_11806 ( .C (clk), .D (new_AGEMA_signal_24529), .Q (new_AGEMA_signal_24530) ) ;
    buf_clk new_AGEMA_reg_buffer_11810 ( .C (clk), .D (new_AGEMA_signal_24533), .Q (new_AGEMA_signal_24534) ) ;
    buf_clk new_AGEMA_reg_buffer_11814 ( .C (clk), .D (new_AGEMA_signal_24537), .Q (new_AGEMA_signal_24538) ) ;
    buf_clk new_AGEMA_reg_buffer_11818 ( .C (clk), .D (new_AGEMA_signal_24541), .Q (new_AGEMA_signal_24542) ) ;
    buf_clk new_AGEMA_reg_buffer_11822 ( .C (clk), .D (new_AGEMA_signal_24545), .Q (new_AGEMA_signal_24546) ) ;
    buf_clk new_AGEMA_reg_buffer_11826 ( .C (clk), .D (new_AGEMA_signal_24549), .Q (new_AGEMA_signal_24550) ) ;
    buf_clk new_AGEMA_reg_buffer_11830 ( .C (clk), .D (new_AGEMA_signal_24553), .Q (new_AGEMA_signal_24554) ) ;
    buf_clk new_AGEMA_reg_buffer_11834 ( .C (clk), .D (new_AGEMA_signal_24557), .Q (new_AGEMA_signal_24558) ) ;
    buf_clk new_AGEMA_reg_buffer_11838 ( .C (clk), .D (new_AGEMA_signal_24561), .Q (new_AGEMA_signal_24562) ) ;
    buf_clk new_AGEMA_reg_buffer_11842 ( .C (clk), .D (new_AGEMA_signal_24565), .Q (new_AGEMA_signal_24566) ) ;
    buf_clk new_AGEMA_reg_buffer_11846 ( .C (clk), .D (new_AGEMA_signal_24569), .Q (new_AGEMA_signal_24570) ) ;
    buf_clk new_AGEMA_reg_buffer_11850 ( .C (clk), .D (new_AGEMA_signal_24573), .Q (new_AGEMA_signal_24574) ) ;
    buf_clk new_AGEMA_reg_buffer_11854 ( .C (clk), .D (new_AGEMA_signal_24577), .Q (new_AGEMA_signal_24578) ) ;
    buf_clk new_AGEMA_reg_buffer_11858 ( .C (clk), .D (new_AGEMA_signal_24581), .Q (new_AGEMA_signal_24582) ) ;
    buf_clk new_AGEMA_reg_buffer_11862 ( .C (clk), .D (new_AGEMA_signal_24585), .Q (new_AGEMA_signal_24586) ) ;
    buf_clk new_AGEMA_reg_buffer_11866 ( .C (clk), .D (new_AGEMA_signal_24589), .Q (new_AGEMA_signal_24590) ) ;
    buf_clk new_AGEMA_reg_buffer_11870 ( .C (clk), .D (new_AGEMA_signal_24593), .Q (new_AGEMA_signal_24594) ) ;
    buf_clk new_AGEMA_reg_buffer_11874 ( .C (clk), .D (new_AGEMA_signal_24597), .Q (new_AGEMA_signal_24598) ) ;
    buf_clk new_AGEMA_reg_buffer_11878 ( .C (clk), .D (new_AGEMA_signal_24601), .Q (new_AGEMA_signal_24602) ) ;
    buf_clk new_AGEMA_reg_buffer_11882 ( .C (clk), .D (new_AGEMA_signal_24605), .Q (new_AGEMA_signal_24606) ) ;
    buf_clk new_AGEMA_reg_buffer_11886 ( .C (clk), .D (new_AGEMA_signal_24609), .Q (new_AGEMA_signal_24610) ) ;
    buf_clk new_AGEMA_reg_buffer_11890 ( .C (clk), .D (new_AGEMA_signal_24613), .Q (new_AGEMA_signal_24614) ) ;
    buf_clk new_AGEMA_reg_buffer_11894 ( .C (clk), .D (new_AGEMA_signal_24617), .Q (new_AGEMA_signal_24618) ) ;
    buf_clk new_AGEMA_reg_buffer_11898 ( .C (clk), .D (new_AGEMA_signal_24621), .Q (new_AGEMA_signal_24622) ) ;
    buf_clk new_AGEMA_reg_buffer_11902 ( .C (clk), .D (new_AGEMA_signal_24625), .Q (new_AGEMA_signal_24626) ) ;
    buf_clk new_AGEMA_reg_buffer_11906 ( .C (clk), .D (new_AGEMA_signal_24629), .Q (new_AGEMA_signal_24630) ) ;
    buf_clk new_AGEMA_reg_buffer_11910 ( .C (clk), .D (new_AGEMA_signal_24633), .Q (new_AGEMA_signal_24634) ) ;
    buf_clk new_AGEMA_reg_buffer_11914 ( .C (clk), .D (new_AGEMA_signal_24637), .Q (new_AGEMA_signal_24638) ) ;
    buf_clk new_AGEMA_reg_buffer_11918 ( .C (clk), .D (new_AGEMA_signal_24641), .Q (new_AGEMA_signal_24642) ) ;
    buf_clk new_AGEMA_reg_buffer_11922 ( .C (clk), .D (new_AGEMA_signal_24645), .Q (new_AGEMA_signal_24646) ) ;
    buf_clk new_AGEMA_reg_buffer_11926 ( .C (clk), .D (new_AGEMA_signal_24649), .Q (new_AGEMA_signal_24650) ) ;
    buf_clk new_AGEMA_reg_buffer_11930 ( .C (clk), .D (new_AGEMA_signal_24653), .Q (new_AGEMA_signal_24654) ) ;
    buf_clk new_AGEMA_reg_buffer_11934 ( .C (clk), .D (new_AGEMA_signal_24657), .Q (new_AGEMA_signal_24658) ) ;
    buf_clk new_AGEMA_reg_buffer_11938 ( .C (clk), .D (new_AGEMA_signal_24661), .Q (new_AGEMA_signal_24662) ) ;
    buf_clk new_AGEMA_reg_buffer_11942 ( .C (clk), .D (new_AGEMA_signal_24665), .Q (new_AGEMA_signal_24666) ) ;
    buf_clk new_AGEMA_reg_buffer_11946 ( .C (clk), .D (new_AGEMA_signal_24669), .Q (new_AGEMA_signal_24670) ) ;
    buf_clk new_AGEMA_reg_buffer_11950 ( .C (clk), .D (new_AGEMA_signal_24673), .Q (new_AGEMA_signal_24674) ) ;
    buf_clk new_AGEMA_reg_buffer_11954 ( .C (clk), .D (new_AGEMA_signal_24677), .Q (new_AGEMA_signal_24678) ) ;
    buf_clk new_AGEMA_reg_buffer_11958 ( .C (clk), .D (new_AGEMA_signal_24681), .Q (new_AGEMA_signal_24682) ) ;
    buf_clk new_AGEMA_reg_buffer_11962 ( .C (clk), .D (new_AGEMA_signal_24685), .Q (new_AGEMA_signal_24686) ) ;
    buf_clk new_AGEMA_reg_buffer_11966 ( .C (clk), .D (new_AGEMA_signal_24689), .Q (new_AGEMA_signal_24690) ) ;
    buf_clk new_AGEMA_reg_buffer_11970 ( .C (clk), .D (new_AGEMA_signal_24693), .Q (new_AGEMA_signal_24694) ) ;
    buf_clk new_AGEMA_reg_buffer_11974 ( .C (clk), .D (new_AGEMA_signal_24697), .Q (new_AGEMA_signal_24698) ) ;
    buf_clk new_AGEMA_reg_buffer_11978 ( .C (clk), .D (new_AGEMA_signal_24701), .Q (new_AGEMA_signal_24702) ) ;
    buf_clk new_AGEMA_reg_buffer_11982 ( .C (clk), .D (new_AGEMA_signal_24705), .Q (new_AGEMA_signal_24706) ) ;
    buf_clk new_AGEMA_reg_buffer_11986 ( .C (clk), .D (new_AGEMA_signal_24709), .Q (new_AGEMA_signal_24710) ) ;
    buf_clk new_AGEMA_reg_buffer_11990 ( .C (clk), .D (new_AGEMA_signal_24713), .Q (new_AGEMA_signal_24714) ) ;
    buf_clk new_AGEMA_reg_buffer_11994 ( .C (clk), .D (new_AGEMA_signal_24717), .Q (new_AGEMA_signal_24718) ) ;
    buf_clk new_AGEMA_reg_buffer_11998 ( .C (clk), .D (new_AGEMA_signal_24721), .Q (new_AGEMA_signal_24722) ) ;
    buf_clk new_AGEMA_reg_buffer_12002 ( .C (clk), .D (new_AGEMA_signal_24725), .Q (new_AGEMA_signal_24726) ) ;
    buf_clk new_AGEMA_reg_buffer_12006 ( .C (clk), .D (new_AGEMA_signal_24729), .Q (new_AGEMA_signal_24730) ) ;
    buf_clk new_AGEMA_reg_buffer_12010 ( .C (clk), .D (new_AGEMA_signal_24733), .Q (new_AGEMA_signal_24734) ) ;
    buf_clk new_AGEMA_reg_buffer_12014 ( .C (clk), .D (new_AGEMA_signal_24737), .Q (new_AGEMA_signal_24738) ) ;
    buf_clk new_AGEMA_reg_buffer_12018 ( .C (clk), .D (new_AGEMA_signal_24741), .Q (new_AGEMA_signal_24742) ) ;
    buf_clk new_AGEMA_reg_buffer_12022 ( .C (clk), .D (new_AGEMA_signal_24745), .Q (new_AGEMA_signal_24746) ) ;
    buf_clk new_AGEMA_reg_buffer_12026 ( .C (clk), .D (new_AGEMA_signal_24749), .Q (new_AGEMA_signal_24750) ) ;
    buf_clk new_AGEMA_reg_buffer_12030 ( .C (clk), .D (new_AGEMA_signal_24753), .Q (new_AGEMA_signal_24754) ) ;
    buf_clk new_AGEMA_reg_buffer_12034 ( .C (clk), .D (new_AGEMA_signal_24757), .Q (new_AGEMA_signal_24758) ) ;
    buf_clk new_AGEMA_reg_buffer_12038 ( .C (clk), .D (new_AGEMA_signal_24761), .Q (new_AGEMA_signal_24762) ) ;
    buf_clk new_AGEMA_reg_buffer_12042 ( .C (clk), .D (new_AGEMA_signal_24765), .Q (new_AGEMA_signal_24766) ) ;
    buf_clk new_AGEMA_reg_buffer_12046 ( .C (clk), .D (new_AGEMA_signal_24769), .Q (new_AGEMA_signal_24770) ) ;
    buf_clk new_AGEMA_reg_buffer_12050 ( .C (clk), .D (new_AGEMA_signal_24773), .Q (new_AGEMA_signal_24774) ) ;
    buf_clk new_AGEMA_reg_buffer_12054 ( .C (clk), .D (new_AGEMA_signal_24777), .Q (new_AGEMA_signal_24778) ) ;
    buf_clk new_AGEMA_reg_buffer_12058 ( .C (clk), .D (new_AGEMA_signal_24781), .Q (new_AGEMA_signal_24782) ) ;
    buf_clk new_AGEMA_reg_buffer_12062 ( .C (clk), .D (new_AGEMA_signal_24785), .Q (new_AGEMA_signal_24786) ) ;
    buf_clk new_AGEMA_reg_buffer_12066 ( .C (clk), .D (new_AGEMA_signal_24789), .Q (new_AGEMA_signal_24790) ) ;
    buf_clk new_AGEMA_reg_buffer_12070 ( .C (clk), .D (new_AGEMA_signal_24793), .Q (new_AGEMA_signal_24794) ) ;
    buf_clk new_AGEMA_reg_buffer_12074 ( .C (clk), .D (new_AGEMA_signal_24797), .Q (new_AGEMA_signal_24798) ) ;
    buf_clk new_AGEMA_reg_buffer_12078 ( .C (clk), .D (new_AGEMA_signal_24801), .Q (new_AGEMA_signal_24802) ) ;
    buf_clk new_AGEMA_reg_buffer_12082 ( .C (clk), .D (new_AGEMA_signal_24805), .Q (new_AGEMA_signal_24806) ) ;
    buf_clk new_AGEMA_reg_buffer_12086 ( .C (clk), .D (new_AGEMA_signal_24809), .Q (new_AGEMA_signal_24810) ) ;
    buf_clk new_AGEMA_reg_buffer_12090 ( .C (clk), .D (new_AGEMA_signal_24813), .Q (new_AGEMA_signal_24814) ) ;
    buf_clk new_AGEMA_reg_buffer_12094 ( .C (clk), .D (new_AGEMA_signal_24817), .Q (new_AGEMA_signal_24818) ) ;
    buf_clk new_AGEMA_reg_buffer_12098 ( .C (clk), .D (new_AGEMA_signal_24821), .Q (new_AGEMA_signal_24822) ) ;
    buf_clk new_AGEMA_reg_buffer_12102 ( .C (clk), .D (new_AGEMA_signal_24825), .Q (new_AGEMA_signal_24826) ) ;
    buf_clk new_AGEMA_reg_buffer_12106 ( .C (clk), .D (new_AGEMA_signal_24829), .Q (new_AGEMA_signal_24830) ) ;
    buf_clk new_AGEMA_reg_buffer_12110 ( .C (clk), .D (new_AGEMA_signal_24833), .Q (new_AGEMA_signal_24834) ) ;
    buf_clk new_AGEMA_reg_buffer_12114 ( .C (clk), .D (new_AGEMA_signal_24837), .Q (new_AGEMA_signal_24838) ) ;
    buf_clk new_AGEMA_reg_buffer_12118 ( .C (clk), .D (new_AGEMA_signal_24841), .Q (new_AGEMA_signal_24842) ) ;
    buf_clk new_AGEMA_reg_buffer_12122 ( .C (clk), .D (new_AGEMA_signal_24845), .Q (new_AGEMA_signal_24846) ) ;
    buf_clk new_AGEMA_reg_buffer_12126 ( .C (clk), .D (new_AGEMA_signal_24849), .Q (new_AGEMA_signal_24850) ) ;
    buf_clk new_AGEMA_reg_buffer_12130 ( .C (clk), .D (new_AGEMA_signal_24853), .Q (new_AGEMA_signal_24854) ) ;
    buf_clk new_AGEMA_reg_buffer_12134 ( .C (clk), .D (new_AGEMA_signal_24857), .Q (new_AGEMA_signal_24858) ) ;
    buf_clk new_AGEMA_reg_buffer_12138 ( .C (clk), .D (new_AGEMA_signal_24861), .Q (new_AGEMA_signal_24862) ) ;
    buf_clk new_AGEMA_reg_buffer_12142 ( .C (clk), .D (new_AGEMA_signal_24865), .Q (new_AGEMA_signal_24866) ) ;
    buf_clk new_AGEMA_reg_buffer_12146 ( .C (clk), .D (new_AGEMA_signal_24869), .Q (new_AGEMA_signal_24870) ) ;
    buf_clk new_AGEMA_reg_buffer_12150 ( .C (clk), .D (new_AGEMA_signal_24873), .Q (new_AGEMA_signal_24874) ) ;
    buf_clk new_AGEMA_reg_buffer_12154 ( .C (clk), .D (new_AGEMA_signal_24877), .Q (new_AGEMA_signal_24878) ) ;
    buf_clk new_AGEMA_reg_buffer_12158 ( .C (clk), .D (new_AGEMA_signal_24881), .Q (new_AGEMA_signal_24882) ) ;
    buf_clk new_AGEMA_reg_buffer_12162 ( .C (clk), .D (new_AGEMA_signal_24885), .Q (new_AGEMA_signal_24886) ) ;
    buf_clk new_AGEMA_reg_buffer_12166 ( .C (clk), .D (new_AGEMA_signal_24889), .Q (new_AGEMA_signal_24890) ) ;
    buf_clk new_AGEMA_reg_buffer_12170 ( .C (clk), .D (new_AGEMA_signal_24893), .Q (new_AGEMA_signal_24894) ) ;
    buf_clk new_AGEMA_reg_buffer_12174 ( .C (clk), .D (new_AGEMA_signal_24897), .Q (new_AGEMA_signal_24898) ) ;
    buf_clk new_AGEMA_reg_buffer_12178 ( .C (clk), .D (new_AGEMA_signal_24901), .Q (new_AGEMA_signal_24902) ) ;
    buf_clk new_AGEMA_reg_buffer_12182 ( .C (clk), .D (new_AGEMA_signal_24905), .Q (new_AGEMA_signal_24906) ) ;
    buf_clk new_AGEMA_reg_buffer_12186 ( .C (clk), .D (new_AGEMA_signal_24909), .Q (new_AGEMA_signal_24910) ) ;
    buf_clk new_AGEMA_reg_buffer_12190 ( .C (clk), .D (new_AGEMA_signal_24913), .Q (new_AGEMA_signal_24914) ) ;
    buf_clk new_AGEMA_reg_buffer_12194 ( .C (clk), .D (new_AGEMA_signal_24917), .Q (new_AGEMA_signal_24918) ) ;
    buf_clk new_AGEMA_reg_buffer_12197 ( .C (clk), .D (new_AGEMA_signal_24920), .Q (new_AGEMA_signal_24921) ) ;
    buf_clk new_AGEMA_reg_buffer_12200 ( .C (clk), .D (new_AGEMA_signal_24923), .Q (new_AGEMA_signal_24924) ) ;
    buf_clk new_AGEMA_reg_buffer_12203 ( .C (clk), .D (new_AGEMA_signal_24926), .Q (new_AGEMA_signal_24927) ) ;
    buf_clk new_AGEMA_reg_buffer_12206 ( .C (clk), .D (new_AGEMA_signal_24929), .Q (new_AGEMA_signal_24930) ) ;
    buf_clk new_AGEMA_reg_buffer_12209 ( .C (clk), .D (new_AGEMA_signal_24932), .Q (new_AGEMA_signal_24933) ) ;
    buf_clk new_AGEMA_reg_buffer_12212 ( .C (clk), .D (new_AGEMA_signal_24935), .Q (new_AGEMA_signal_24936) ) ;
    buf_clk new_AGEMA_reg_buffer_12215 ( .C (clk), .D (new_AGEMA_signal_24938), .Q (new_AGEMA_signal_24939) ) ;
    buf_clk new_AGEMA_reg_buffer_12218 ( .C (clk), .D (new_AGEMA_signal_24941), .Q (new_AGEMA_signal_24942) ) ;
    buf_clk new_AGEMA_reg_buffer_12221 ( .C (clk), .D (new_AGEMA_signal_24944), .Q (new_AGEMA_signal_24945) ) ;
    buf_clk new_AGEMA_reg_buffer_12224 ( .C (clk), .D (new_AGEMA_signal_24947), .Q (new_AGEMA_signal_24948) ) ;
    buf_clk new_AGEMA_reg_buffer_12227 ( .C (clk), .D (new_AGEMA_signal_24950), .Q (new_AGEMA_signal_24951) ) ;
    buf_clk new_AGEMA_reg_buffer_12230 ( .C (clk), .D (new_AGEMA_signal_24953), .Q (new_AGEMA_signal_24954) ) ;
    buf_clk new_AGEMA_reg_buffer_12233 ( .C (clk), .D (new_AGEMA_signal_24956), .Q (new_AGEMA_signal_24957) ) ;
    buf_clk new_AGEMA_reg_buffer_12236 ( .C (clk), .D (new_AGEMA_signal_24959), .Q (new_AGEMA_signal_24960) ) ;
    buf_clk new_AGEMA_reg_buffer_12239 ( .C (clk), .D (new_AGEMA_signal_24962), .Q (new_AGEMA_signal_24963) ) ;
    buf_clk new_AGEMA_reg_buffer_12242 ( .C (clk), .D (new_AGEMA_signal_24965), .Q (new_AGEMA_signal_24966) ) ;
    buf_clk new_AGEMA_reg_buffer_12245 ( .C (clk), .D (new_AGEMA_signal_24968), .Q (new_AGEMA_signal_24969) ) ;
    buf_clk new_AGEMA_reg_buffer_12248 ( .C (clk), .D (new_AGEMA_signal_24971), .Q (new_AGEMA_signal_24972) ) ;
    buf_clk new_AGEMA_reg_buffer_12251 ( .C (clk), .D (new_AGEMA_signal_24974), .Q (new_AGEMA_signal_24975) ) ;
    buf_clk new_AGEMA_reg_buffer_12254 ( .C (clk), .D (new_AGEMA_signal_24977), .Q (new_AGEMA_signal_24978) ) ;
    buf_clk new_AGEMA_reg_buffer_12257 ( .C (clk), .D (new_AGEMA_signal_24980), .Q (new_AGEMA_signal_24981) ) ;
    buf_clk new_AGEMA_reg_buffer_12260 ( .C (clk), .D (new_AGEMA_signal_24983), .Q (new_AGEMA_signal_24984) ) ;
    buf_clk new_AGEMA_reg_buffer_12263 ( .C (clk), .D (new_AGEMA_signal_24986), .Q (new_AGEMA_signal_24987) ) ;
    buf_clk new_AGEMA_reg_buffer_12266 ( .C (clk), .D (new_AGEMA_signal_24989), .Q (new_AGEMA_signal_24990) ) ;
    buf_clk new_AGEMA_reg_buffer_12269 ( .C (clk), .D (new_AGEMA_signal_24992), .Q (new_AGEMA_signal_24993) ) ;
    buf_clk new_AGEMA_reg_buffer_12272 ( .C (clk), .D (new_AGEMA_signal_24995), .Q (new_AGEMA_signal_24996) ) ;
    buf_clk new_AGEMA_reg_buffer_12275 ( .C (clk), .D (new_AGEMA_signal_24998), .Q (new_AGEMA_signal_24999) ) ;
    buf_clk new_AGEMA_reg_buffer_12278 ( .C (clk), .D (new_AGEMA_signal_25001), .Q (new_AGEMA_signal_25002) ) ;
    buf_clk new_AGEMA_reg_buffer_12281 ( .C (clk), .D (new_AGEMA_signal_25004), .Q (new_AGEMA_signal_25005) ) ;
    buf_clk new_AGEMA_reg_buffer_12284 ( .C (clk), .D (new_AGEMA_signal_25007), .Q (new_AGEMA_signal_25008) ) ;
    buf_clk new_AGEMA_reg_buffer_12287 ( .C (clk), .D (new_AGEMA_signal_25010), .Q (new_AGEMA_signal_25011) ) ;
    buf_clk new_AGEMA_reg_buffer_12290 ( .C (clk), .D (new_AGEMA_signal_25013), .Q (new_AGEMA_signal_25014) ) ;
    buf_clk new_AGEMA_reg_buffer_12293 ( .C (clk), .D (new_AGEMA_signal_25016), .Q (new_AGEMA_signal_25017) ) ;
    buf_clk new_AGEMA_reg_buffer_12296 ( .C (clk), .D (new_AGEMA_signal_25019), .Q (new_AGEMA_signal_25020) ) ;
    buf_clk new_AGEMA_reg_buffer_12299 ( .C (clk), .D (new_AGEMA_signal_25022), .Q (new_AGEMA_signal_25023) ) ;
    buf_clk new_AGEMA_reg_buffer_12302 ( .C (clk), .D (new_AGEMA_signal_25025), .Q (new_AGEMA_signal_25026) ) ;
    buf_clk new_AGEMA_reg_buffer_12305 ( .C (clk), .D (new_AGEMA_signal_25028), .Q (new_AGEMA_signal_25029) ) ;
    buf_clk new_AGEMA_reg_buffer_12308 ( .C (clk), .D (new_AGEMA_signal_25031), .Q (new_AGEMA_signal_25032) ) ;
    buf_clk new_AGEMA_reg_buffer_12311 ( .C (clk), .D (new_AGEMA_signal_25034), .Q (new_AGEMA_signal_25035) ) ;
    buf_clk new_AGEMA_reg_buffer_12314 ( .C (clk), .D (new_AGEMA_signal_25037), .Q (new_AGEMA_signal_25038) ) ;
    buf_clk new_AGEMA_reg_buffer_12317 ( .C (clk), .D (new_AGEMA_signal_25040), .Q (new_AGEMA_signal_25041) ) ;
    buf_clk new_AGEMA_reg_buffer_12320 ( .C (clk), .D (new_AGEMA_signal_25043), .Q (new_AGEMA_signal_25044) ) ;
    buf_clk new_AGEMA_reg_buffer_12323 ( .C (clk), .D (new_AGEMA_signal_25046), .Q (new_AGEMA_signal_25047) ) ;
    buf_clk new_AGEMA_reg_buffer_12326 ( .C (clk), .D (new_AGEMA_signal_25049), .Q (new_AGEMA_signal_25050) ) ;
    buf_clk new_AGEMA_reg_buffer_12329 ( .C (clk), .D (new_AGEMA_signal_25052), .Q (new_AGEMA_signal_25053) ) ;
    buf_clk new_AGEMA_reg_buffer_12332 ( .C (clk), .D (new_AGEMA_signal_25055), .Q (new_AGEMA_signal_25056) ) ;
    buf_clk new_AGEMA_reg_buffer_12335 ( .C (clk), .D (new_AGEMA_signal_25058), .Q (new_AGEMA_signal_25059) ) ;
    buf_clk new_AGEMA_reg_buffer_12338 ( .C (clk), .D (new_AGEMA_signal_25061), .Q (new_AGEMA_signal_25062) ) ;
    buf_clk new_AGEMA_reg_buffer_12341 ( .C (clk), .D (new_AGEMA_signal_25064), .Q (new_AGEMA_signal_25065) ) ;
    buf_clk new_AGEMA_reg_buffer_12344 ( .C (clk), .D (new_AGEMA_signal_25067), .Q (new_AGEMA_signal_25068) ) ;
    buf_clk new_AGEMA_reg_buffer_12347 ( .C (clk), .D (new_AGEMA_signal_25070), .Q (new_AGEMA_signal_25071) ) ;
    buf_clk new_AGEMA_reg_buffer_12350 ( .C (clk), .D (new_AGEMA_signal_25073), .Q (new_AGEMA_signal_25074) ) ;
    buf_clk new_AGEMA_reg_buffer_12353 ( .C (clk), .D (new_AGEMA_signal_25076), .Q (new_AGEMA_signal_25077) ) ;
    buf_clk new_AGEMA_reg_buffer_12356 ( .C (clk), .D (new_AGEMA_signal_25079), .Q (new_AGEMA_signal_25080) ) ;
    buf_clk new_AGEMA_reg_buffer_12359 ( .C (clk), .D (new_AGEMA_signal_25082), .Q (new_AGEMA_signal_25083) ) ;
    buf_clk new_AGEMA_reg_buffer_12362 ( .C (clk), .D (new_AGEMA_signal_25085), .Q (new_AGEMA_signal_25086) ) ;
    buf_clk new_AGEMA_reg_buffer_12365 ( .C (clk), .D (new_AGEMA_signal_25088), .Q (new_AGEMA_signal_25089) ) ;
    buf_clk new_AGEMA_reg_buffer_12368 ( .C (clk), .D (new_AGEMA_signal_25091), .Q (new_AGEMA_signal_25092) ) ;
    buf_clk new_AGEMA_reg_buffer_12371 ( .C (clk), .D (new_AGEMA_signal_25094), .Q (new_AGEMA_signal_25095) ) ;
    buf_clk new_AGEMA_reg_buffer_12374 ( .C (clk), .D (new_AGEMA_signal_25097), .Q (new_AGEMA_signal_25098) ) ;
    buf_clk new_AGEMA_reg_buffer_12377 ( .C (clk), .D (new_AGEMA_signal_25100), .Q (new_AGEMA_signal_25101) ) ;
    buf_clk new_AGEMA_reg_buffer_12380 ( .C (clk), .D (new_AGEMA_signal_25103), .Q (new_AGEMA_signal_25104) ) ;
    buf_clk new_AGEMA_reg_buffer_12383 ( .C (clk), .D (new_AGEMA_signal_25106), .Q (new_AGEMA_signal_25107) ) ;
    buf_clk new_AGEMA_reg_buffer_12386 ( .C (clk), .D (new_AGEMA_signal_25109), .Q (new_AGEMA_signal_25110) ) ;
    buf_clk new_AGEMA_reg_buffer_12389 ( .C (clk), .D (new_AGEMA_signal_25112), .Q (new_AGEMA_signal_25113) ) ;
    buf_clk new_AGEMA_reg_buffer_12392 ( .C (clk), .D (new_AGEMA_signal_25115), .Q (new_AGEMA_signal_25116) ) ;
    buf_clk new_AGEMA_reg_buffer_12395 ( .C (clk), .D (new_AGEMA_signal_25118), .Q (new_AGEMA_signal_25119) ) ;
    buf_clk new_AGEMA_reg_buffer_12398 ( .C (clk), .D (new_AGEMA_signal_25121), .Q (new_AGEMA_signal_25122) ) ;
    buf_clk new_AGEMA_reg_buffer_12401 ( .C (clk), .D (new_AGEMA_signal_25124), .Q (new_AGEMA_signal_25125) ) ;
    buf_clk new_AGEMA_reg_buffer_12404 ( .C (clk), .D (new_AGEMA_signal_25127), .Q (new_AGEMA_signal_25128) ) ;
    buf_clk new_AGEMA_reg_buffer_12407 ( .C (clk), .D (new_AGEMA_signal_25130), .Q (new_AGEMA_signal_25131) ) ;
    buf_clk new_AGEMA_reg_buffer_12410 ( .C (clk), .D (new_AGEMA_signal_25133), .Q (new_AGEMA_signal_25134) ) ;
    buf_clk new_AGEMA_reg_buffer_12413 ( .C (clk), .D (new_AGEMA_signal_25136), .Q (new_AGEMA_signal_25137) ) ;
    buf_clk new_AGEMA_reg_buffer_12416 ( .C (clk), .D (new_AGEMA_signal_25139), .Q (new_AGEMA_signal_25140) ) ;
    buf_clk new_AGEMA_reg_buffer_12419 ( .C (clk), .D (new_AGEMA_signal_25142), .Q (new_AGEMA_signal_25143) ) ;
    buf_clk new_AGEMA_reg_buffer_12422 ( .C (clk), .D (new_AGEMA_signal_25145), .Q (new_AGEMA_signal_25146) ) ;
    buf_clk new_AGEMA_reg_buffer_12425 ( .C (clk), .D (new_AGEMA_signal_25148), .Q (new_AGEMA_signal_25149) ) ;
    buf_clk new_AGEMA_reg_buffer_12428 ( .C (clk), .D (new_AGEMA_signal_25151), .Q (new_AGEMA_signal_25152) ) ;
    buf_clk new_AGEMA_reg_buffer_12431 ( .C (clk), .D (new_AGEMA_signal_25154), .Q (new_AGEMA_signal_25155) ) ;
    buf_clk new_AGEMA_reg_buffer_12434 ( .C (clk), .D (new_AGEMA_signal_25157), .Q (new_AGEMA_signal_25158) ) ;
    buf_clk new_AGEMA_reg_buffer_12437 ( .C (clk), .D (new_AGEMA_signal_25160), .Q (new_AGEMA_signal_25161) ) ;
    buf_clk new_AGEMA_reg_buffer_12440 ( .C (clk), .D (new_AGEMA_signal_25163), .Q (new_AGEMA_signal_25164) ) ;
    buf_clk new_AGEMA_reg_buffer_12443 ( .C (clk), .D (new_AGEMA_signal_25166), .Q (new_AGEMA_signal_25167) ) ;
    buf_clk new_AGEMA_reg_buffer_12446 ( .C (clk), .D (new_AGEMA_signal_25169), .Q (new_AGEMA_signal_25170) ) ;
    buf_clk new_AGEMA_reg_buffer_12449 ( .C (clk), .D (new_AGEMA_signal_25172), .Q (new_AGEMA_signal_25173) ) ;
    buf_clk new_AGEMA_reg_buffer_12452 ( .C (clk), .D (new_AGEMA_signal_25175), .Q (new_AGEMA_signal_25176) ) ;
    buf_clk new_AGEMA_reg_buffer_12455 ( .C (clk), .D (new_AGEMA_signal_25178), .Q (new_AGEMA_signal_25179) ) ;
    buf_clk new_AGEMA_reg_buffer_12458 ( .C (clk), .D (new_AGEMA_signal_25181), .Q (new_AGEMA_signal_25182) ) ;
    buf_clk new_AGEMA_reg_buffer_12461 ( .C (clk), .D (new_AGEMA_signal_25184), .Q (new_AGEMA_signal_25185) ) ;
    buf_clk new_AGEMA_reg_buffer_12464 ( .C (clk), .D (new_AGEMA_signal_25187), .Q (new_AGEMA_signal_25188) ) ;
    buf_clk new_AGEMA_reg_buffer_12467 ( .C (clk), .D (new_AGEMA_signal_25190), .Q (new_AGEMA_signal_25191) ) ;
    buf_clk new_AGEMA_reg_buffer_12470 ( .C (clk), .D (new_AGEMA_signal_25193), .Q (new_AGEMA_signal_25194) ) ;
    buf_clk new_AGEMA_reg_buffer_12473 ( .C (clk), .D (new_AGEMA_signal_25196), .Q (new_AGEMA_signal_25197) ) ;
    buf_clk new_AGEMA_reg_buffer_12476 ( .C (clk), .D (new_AGEMA_signal_25199), .Q (new_AGEMA_signal_25200) ) ;
    buf_clk new_AGEMA_reg_buffer_12479 ( .C (clk), .D (new_AGEMA_signal_25202), .Q (new_AGEMA_signal_25203) ) ;
    buf_clk new_AGEMA_reg_buffer_12482 ( .C (clk), .D (new_AGEMA_signal_25205), .Q (new_AGEMA_signal_25206) ) ;
    buf_clk new_AGEMA_reg_buffer_12485 ( .C (clk), .D (new_AGEMA_signal_25208), .Q (new_AGEMA_signal_25209) ) ;
    buf_clk new_AGEMA_reg_buffer_12488 ( .C (clk), .D (new_AGEMA_signal_25211), .Q (new_AGEMA_signal_25212) ) ;
    buf_clk new_AGEMA_reg_buffer_12491 ( .C (clk), .D (new_AGEMA_signal_25214), .Q (new_AGEMA_signal_25215) ) ;
    buf_clk new_AGEMA_reg_buffer_12494 ( .C (clk), .D (new_AGEMA_signal_25217), .Q (new_AGEMA_signal_25218) ) ;
    buf_clk new_AGEMA_reg_buffer_12497 ( .C (clk), .D (new_AGEMA_signal_25220), .Q (new_AGEMA_signal_25221) ) ;
    buf_clk new_AGEMA_reg_buffer_12500 ( .C (clk), .D (new_AGEMA_signal_25223), .Q (new_AGEMA_signal_25224) ) ;
    buf_clk new_AGEMA_reg_buffer_12503 ( .C (clk), .D (new_AGEMA_signal_25226), .Q (new_AGEMA_signal_25227) ) ;
    buf_clk new_AGEMA_reg_buffer_12506 ( .C (clk), .D (new_AGEMA_signal_25229), .Q (new_AGEMA_signal_25230) ) ;
    buf_clk new_AGEMA_reg_buffer_12509 ( .C (clk), .D (new_AGEMA_signal_25232), .Q (new_AGEMA_signal_25233) ) ;
    buf_clk new_AGEMA_reg_buffer_12512 ( .C (clk), .D (new_AGEMA_signal_25235), .Q (new_AGEMA_signal_25236) ) ;
    buf_clk new_AGEMA_reg_buffer_12515 ( .C (clk), .D (new_AGEMA_signal_25238), .Q (new_AGEMA_signal_25239) ) ;
    buf_clk new_AGEMA_reg_buffer_12518 ( .C (clk), .D (new_AGEMA_signal_25241), .Q (new_AGEMA_signal_25242) ) ;
    buf_clk new_AGEMA_reg_buffer_12521 ( .C (clk), .D (new_AGEMA_signal_25244), .Q (new_AGEMA_signal_25245) ) ;
    buf_clk new_AGEMA_reg_buffer_12524 ( .C (clk), .D (new_AGEMA_signal_25247), .Q (new_AGEMA_signal_25248) ) ;
    buf_clk new_AGEMA_reg_buffer_12527 ( .C (clk), .D (new_AGEMA_signal_25250), .Q (new_AGEMA_signal_25251) ) ;
    buf_clk new_AGEMA_reg_buffer_12530 ( .C (clk), .D (new_AGEMA_signal_25253), .Q (new_AGEMA_signal_25254) ) ;
    buf_clk new_AGEMA_reg_buffer_12533 ( .C (clk), .D (new_AGEMA_signal_25256), .Q (new_AGEMA_signal_25257) ) ;
    buf_clk new_AGEMA_reg_buffer_12536 ( .C (clk), .D (new_AGEMA_signal_25259), .Q (new_AGEMA_signal_25260) ) ;
    buf_clk new_AGEMA_reg_buffer_12539 ( .C (clk), .D (new_AGEMA_signal_25262), .Q (new_AGEMA_signal_25263) ) ;
    buf_clk new_AGEMA_reg_buffer_12542 ( .C (clk), .D (new_AGEMA_signal_25265), .Q (new_AGEMA_signal_25266) ) ;
    buf_clk new_AGEMA_reg_buffer_12545 ( .C (clk), .D (new_AGEMA_signal_25268), .Q (new_AGEMA_signal_25269) ) ;
    buf_clk new_AGEMA_reg_buffer_12548 ( .C (clk), .D (new_AGEMA_signal_25271), .Q (new_AGEMA_signal_25272) ) ;
    buf_clk new_AGEMA_reg_buffer_12551 ( .C (clk), .D (new_AGEMA_signal_25274), .Q (new_AGEMA_signal_25275) ) ;
    buf_clk new_AGEMA_reg_buffer_12554 ( .C (clk), .D (new_AGEMA_signal_25277), .Q (new_AGEMA_signal_25278) ) ;
    buf_clk new_AGEMA_reg_buffer_12557 ( .C (clk), .D (new_AGEMA_signal_25280), .Q (new_AGEMA_signal_25281) ) ;
    buf_clk new_AGEMA_reg_buffer_12560 ( .C (clk), .D (new_AGEMA_signal_25283), .Q (new_AGEMA_signal_25284) ) ;
    buf_clk new_AGEMA_reg_buffer_12563 ( .C (clk), .D (new_AGEMA_signal_25286), .Q (new_AGEMA_signal_25287) ) ;
    buf_clk new_AGEMA_reg_buffer_12566 ( .C (clk), .D (new_AGEMA_signal_25289), .Q (new_AGEMA_signal_25290) ) ;
    buf_clk new_AGEMA_reg_buffer_12569 ( .C (clk), .D (new_AGEMA_signal_25292), .Q (new_AGEMA_signal_25293) ) ;
    buf_clk new_AGEMA_reg_buffer_12572 ( .C (clk), .D (new_AGEMA_signal_25295), .Q (new_AGEMA_signal_25296) ) ;
    buf_clk new_AGEMA_reg_buffer_12575 ( .C (clk), .D (new_AGEMA_signal_25298), .Q (new_AGEMA_signal_25299) ) ;
    buf_clk new_AGEMA_reg_buffer_12578 ( .C (clk), .D (new_AGEMA_signal_25301), .Q (new_AGEMA_signal_25302) ) ;
    buf_clk new_AGEMA_reg_buffer_12581 ( .C (clk), .D (new_AGEMA_signal_25304), .Q (new_AGEMA_signal_25305) ) ;
    buf_clk new_AGEMA_reg_buffer_12584 ( .C (clk), .D (new_AGEMA_signal_25307), .Q (new_AGEMA_signal_25308) ) ;
    buf_clk new_AGEMA_reg_buffer_12587 ( .C (clk), .D (new_AGEMA_signal_25310), .Q (new_AGEMA_signal_25311) ) ;
    buf_clk new_AGEMA_reg_buffer_12590 ( .C (clk), .D (new_AGEMA_signal_25313), .Q (new_AGEMA_signal_25314) ) ;
    buf_clk new_AGEMA_reg_buffer_12593 ( .C (clk), .D (new_AGEMA_signal_25316), .Q (new_AGEMA_signal_25317) ) ;
    buf_clk new_AGEMA_reg_buffer_12596 ( .C (clk), .D (new_AGEMA_signal_25319), .Q (new_AGEMA_signal_25320) ) ;
    buf_clk new_AGEMA_reg_buffer_12599 ( .C (clk), .D (new_AGEMA_signal_25322), .Q (new_AGEMA_signal_25323) ) ;
    buf_clk new_AGEMA_reg_buffer_12602 ( .C (clk), .D (new_AGEMA_signal_25325), .Q (new_AGEMA_signal_25326) ) ;
    buf_clk new_AGEMA_reg_buffer_12605 ( .C (clk), .D (new_AGEMA_signal_25328), .Q (new_AGEMA_signal_25329) ) ;
    buf_clk new_AGEMA_reg_buffer_12608 ( .C (clk), .D (new_AGEMA_signal_25331), .Q (new_AGEMA_signal_25332) ) ;
    buf_clk new_AGEMA_reg_buffer_12611 ( .C (clk), .D (new_AGEMA_signal_25334), .Q (new_AGEMA_signal_25335) ) ;
    buf_clk new_AGEMA_reg_buffer_12614 ( .C (clk), .D (new_AGEMA_signal_25337), .Q (new_AGEMA_signal_25338) ) ;
    buf_clk new_AGEMA_reg_buffer_12617 ( .C (clk), .D (new_AGEMA_signal_25340), .Q (new_AGEMA_signal_25341) ) ;
    buf_clk new_AGEMA_reg_buffer_12620 ( .C (clk), .D (new_AGEMA_signal_25343), .Q (new_AGEMA_signal_25344) ) ;
    buf_clk new_AGEMA_reg_buffer_12623 ( .C (clk), .D (new_AGEMA_signal_25346), .Q (new_AGEMA_signal_25347) ) ;
    buf_clk new_AGEMA_reg_buffer_12626 ( .C (clk), .D (new_AGEMA_signal_25349), .Q (new_AGEMA_signal_25350) ) ;
    buf_clk new_AGEMA_reg_buffer_12629 ( .C (clk), .D (new_AGEMA_signal_25352), .Q (new_AGEMA_signal_25353) ) ;
    buf_clk new_AGEMA_reg_buffer_12632 ( .C (clk), .D (new_AGEMA_signal_25355), .Q (new_AGEMA_signal_25356) ) ;
    buf_clk new_AGEMA_reg_buffer_12635 ( .C (clk), .D (new_AGEMA_signal_25358), .Q (new_AGEMA_signal_25359) ) ;
    buf_clk new_AGEMA_reg_buffer_12638 ( .C (clk), .D (new_AGEMA_signal_25361), .Q (new_AGEMA_signal_25362) ) ;
    buf_clk new_AGEMA_reg_buffer_12641 ( .C (clk), .D (new_AGEMA_signal_25364), .Q (new_AGEMA_signal_25365) ) ;
    buf_clk new_AGEMA_reg_buffer_12644 ( .C (clk), .D (new_AGEMA_signal_25367), .Q (new_AGEMA_signal_25368) ) ;
    buf_clk new_AGEMA_reg_buffer_12647 ( .C (clk), .D (new_AGEMA_signal_25370), .Q (new_AGEMA_signal_25371) ) ;
    buf_clk new_AGEMA_reg_buffer_12650 ( .C (clk), .D (new_AGEMA_signal_25373), .Q (new_AGEMA_signal_25374) ) ;
    buf_clk new_AGEMA_reg_buffer_12653 ( .C (clk), .D (new_AGEMA_signal_25376), .Q (new_AGEMA_signal_25377) ) ;
    buf_clk new_AGEMA_reg_buffer_12656 ( .C (clk), .D (new_AGEMA_signal_25379), .Q (new_AGEMA_signal_25380) ) ;
    buf_clk new_AGEMA_reg_buffer_12659 ( .C (clk), .D (new_AGEMA_signal_25382), .Q (new_AGEMA_signal_25383) ) ;
    buf_clk new_AGEMA_reg_buffer_12662 ( .C (clk), .D (new_AGEMA_signal_25385), .Q (new_AGEMA_signal_25386) ) ;
    buf_clk new_AGEMA_reg_buffer_12665 ( .C (clk), .D (new_AGEMA_signal_25388), .Q (new_AGEMA_signal_25389) ) ;
    buf_clk new_AGEMA_reg_buffer_12668 ( .C (clk), .D (new_AGEMA_signal_25391), .Q (new_AGEMA_signal_25392) ) ;
    buf_clk new_AGEMA_reg_buffer_12671 ( .C (clk), .D (new_AGEMA_signal_25394), .Q (new_AGEMA_signal_25395) ) ;
    buf_clk new_AGEMA_reg_buffer_12674 ( .C (clk), .D (new_AGEMA_signal_25397), .Q (new_AGEMA_signal_25398) ) ;
    buf_clk new_AGEMA_reg_buffer_12677 ( .C (clk), .D (new_AGEMA_signal_25400), .Q (new_AGEMA_signal_25401) ) ;
    buf_clk new_AGEMA_reg_buffer_12680 ( .C (clk), .D (new_AGEMA_signal_25403), .Q (new_AGEMA_signal_25404) ) ;
    buf_clk new_AGEMA_reg_buffer_12683 ( .C (clk), .D (new_AGEMA_signal_25406), .Q (new_AGEMA_signal_25407) ) ;
    buf_clk new_AGEMA_reg_buffer_12686 ( .C (clk), .D (new_AGEMA_signal_25409), .Q (new_AGEMA_signal_25410) ) ;
    buf_clk new_AGEMA_reg_buffer_12689 ( .C (clk), .D (new_AGEMA_signal_25412), .Q (new_AGEMA_signal_25413) ) ;
    buf_clk new_AGEMA_reg_buffer_12692 ( .C (clk), .D (new_AGEMA_signal_25415), .Q (new_AGEMA_signal_25416) ) ;
    buf_clk new_AGEMA_reg_buffer_12695 ( .C (clk), .D (new_AGEMA_signal_25418), .Q (new_AGEMA_signal_25419) ) ;
    buf_clk new_AGEMA_reg_buffer_12698 ( .C (clk), .D (new_AGEMA_signal_25421), .Q (new_AGEMA_signal_25422) ) ;
    buf_clk new_AGEMA_reg_buffer_12701 ( .C (clk), .D (new_AGEMA_signal_25424), .Q (new_AGEMA_signal_25425) ) ;
    buf_clk new_AGEMA_reg_buffer_12704 ( .C (clk), .D (new_AGEMA_signal_25427), .Q (new_AGEMA_signal_25428) ) ;
    buf_clk new_AGEMA_reg_buffer_12707 ( .C (clk), .D (new_AGEMA_signal_25430), .Q (new_AGEMA_signal_25431) ) ;
    buf_clk new_AGEMA_reg_buffer_12710 ( .C (clk), .D (new_AGEMA_signal_25433), .Q (new_AGEMA_signal_25434) ) ;
    buf_clk new_AGEMA_reg_buffer_12713 ( .C (clk), .D (new_AGEMA_signal_25436), .Q (new_AGEMA_signal_25437) ) ;
    buf_clk new_AGEMA_reg_buffer_12716 ( .C (clk), .D (new_AGEMA_signal_25439), .Q (new_AGEMA_signal_25440) ) ;
    buf_clk new_AGEMA_reg_buffer_12719 ( .C (clk), .D (new_AGEMA_signal_25442), .Q (new_AGEMA_signal_25443) ) ;
    buf_clk new_AGEMA_reg_buffer_12722 ( .C (clk), .D (new_AGEMA_signal_25445), .Q (new_AGEMA_signal_25446) ) ;
    buf_clk new_AGEMA_reg_buffer_12725 ( .C (clk), .D (new_AGEMA_signal_25448), .Q (new_AGEMA_signal_25449) ) ;
    buf_clk new_AGEMA_reg_buffer_12728 ( .C (clk), .D (new_AGEMA_signal_25451), .Q (new_AGEMA_signal_25452) ) ;
    buf_clk new_AGEMA_reg_buffer_12731 ( .C (clk), .D (new_AGEMA_signal_25454), .Q (new_AGEMA_signal_25455) ) ;
    buf_clk new_AGEMA_reg_buffer_12734 ( .C (clk), .D (new_AGEMA_signal_25457), .Q (new_AGEMA_signal_25458) ) ;
    buf_clk new_AGEMA_reg_buffer_12737 ( .C (clk), .D (new_AGEMA_signal_25460), .Q (new_AGEMA_signal_25461) ) ;
    buf_clk new_AGEMA_reg_buffer_12740 ( .C (clk), .D (new_AGEMA_signal_25463), .Q (new_AGEMA_signal_25464) ) ;
    buf_clk new_AGEMA_reg_buffer_12743 ( .C (clk), .D (new_AGEMA_signal_25466), .Q (new_AGEMA_signal_25467) ) ;
    buf_clk new_AGEMA_reg_buffer_12746 ( .C (clk), .D (new_AGEMA_signal_25469), .Q (new_AGEMA_signal_25470) ) ;
    buf_clk new_AGEMA_reg_buffer_12749 ( .C (clk), .D (new_AGEMA_signal_25472), .Q (new_AGEMA_signal_25473) ) ;
    buf_clk new_AGEMA_reg_buffer_12752 ( .C (clk), .D (new_AGEMA_signal_25475), .Q (new_AGEMA_signal_25476) ) ;
    buf_clk new_AGEMA_reg_buffer_12755 ( .C (clk), .D (new_AGEMA_signal_25478), .Q (new_AGEMA_signal_25479) ) ;
    buf_clk new_AGEMA_reg_buffer_12758 ( .C (clk), .D (new_AGEMA_signal_25481), .Q (new_AGEMA_signal_25482) ) ;
    buf_clk new_AGEMA_reg_buffer_12761 ( .C (clk), .D (new_AGEMA_signal_25484), .Q (new_AGEMA_signal_25485) ) ;
    buf_clk new_AGEMA_reg_buffer_12764 ( .C (clk), .D (new_AGEMA_signal_25487), .Q (new_AGEMA_signal_25488) ) ;
    buf_clk new_AGEMA_reg_buffer_12767 ( .C (clk), .D (new_AGEMA_signal_25490), .Q (new_AGEMA_signal_25491) ) ;
    buf_clk new_AGEMA_reg_buffer_12770 ( .C (clk), .D (new_AGEMA_signal_25493), .Q (new_AGEMA_signal_25494) ) ;
    buf_clk new_AGEMA_reg_buffer_12773 ( .C (clk), .D (new_AGEMA_signal_25496), .Q (new_AGEMA_signal_25497) ) ;
    buf_clk new_AGEMA_reg_buffer_12776 ( .C (clk), .D (new_AGEMA_signal_25499), .Q (new_AGEMA_signal_25500) ) ;
    buf_clk new_AGEMA_reg_buffer_12779 ( .C (clk), .D (new_AGEMA_signal_25502), .Q (new_AGEMA_signal_25503) ) ;
    buf_clk new_AGEMA_reg_buffer_12782 ( .C (clk), .D (new_AGEMA_signal_25505), .Q (new_AGEMA_signal_25506) ) ;
    buf_clk new_AGEMA_reg_buffer_12785 ( .C (clk), .D (new_AGEMA_signal_25508), .Q (new_AGEMA_signal_25509) ) ;
    buf_clk new_AGEMA_reg_buffer_12788 ( .C (clk), .D (new_AGEMA_signal_25511), .Q (new_AGEMA_signal_25512) ) ;
    buf_clk new_AGEMA_reg_buffer_12791 ( .C (clk), .D (new_AGEMA_signal_25514), .Q (new_AGEMA_signal_25515) ) ;
    buf_clk new_AGEMA_reg_buffer_12794 ( .C (clk), .D (new_AGEMA_signal_25517), .Q (new_AGEMA_signal_25518) ) ;
    buf_clk new_AGEMA_reg_buffer_12797 ( .C (clk), .D (new_AGEMA_signal_25520), .Q (new_AGEMA_signal_25521) ) ;
    buf_clk new_AGEMA_reg_buffer_12800 ( .C (clk), .D (new_AGEMA_signal_25523), .Q (new_AGEMA_signal_25524) ) ;
    buf_clk new_AGEMA_reg_buffer_12803 ( .C (clk), .D (new_AGEMA_signal_25526), .Q (new_AGEMA_signal_25527) ) ;
    buf_clk new_AGEMA_reg_buffer_12806 ( .C (clk), .D (new_AGEMA_signal_25529), .Q (new_AGEMA_signal_25530) ) ;
    buf_clk new_AGEMA_reg_buffer_12810 ( .C (clk), .D (new_AGEMA_signal_25533), .Q (new_AGEMA_signal_25534) ) ;
    buf_clk new_AGEMA_reg_buffer_12814 ( .C (clk), .D (new_AGEMA_signal_25537), .Q (new_AGEMA_signal_25538) ) ;
    buf_clk new_AGEMA_reg_buffer_12818 ( .C (clk), .D (new_AGEMA_signal_25541), .Q (new_AGEMA_signal_25542) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_17181, new_AGEMA_signal_17180, new_AGEMA_signal_17179}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_17184, new_AGEMA_signal_17183, new_AGEMA_signal_17182}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_17181, new_AGEMA_signal_17180, new_AGEMA_signal_17179}), .b ({new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_17184, new_AGEMA_signal_17183, new_AGEMA_signal_17182}), .b ({new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_17415, new_AGEMA_signal_17414, new_AGEMA_signal_17413}), .b ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_17418, new_AGEMA_signal_17417, new_AGEMA_signal_17416}), .c ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_17421, new_AGEMA_signal_17420, new_AGEMA_signal_17419}), .b ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_17424, new_AGEMA_signal_17423, new_AGEMA_signal_17422}), .c ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_17193, new_AGEMA_signal_17192, new_AGEMA_signal_17191}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_17196, new_AGEMA_signal_17195, new_AGEMA_signal_17194}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_17193, new_AGEMA_signal_17192, new_AGEMA_signal_17191}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_17196, new_AGEMA_signal_17195, new_AGEMA_signal_17194}), .b ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_17427, new_AGEMA_signal_17426, new_AGEMA_signal_17425}), .b ({new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_17430, new_AGEMA_signal_17429, new_AGEMA_signal_17428}), .c ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_17433, new_AGEMA_signal_17432, new_AGEMA_signal_17431}), .b ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_17436, new_AGEMA_signal_17435, new_AGEMA_signal_17434}), .c ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_17205, new_AGEMA_signal_17204, new_AGEMA_signal_17203}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_17208, new_AGEMA_signal_17207, new_AGEMA_signal_17206}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_17205, new_AGEMA_signal_17204, new_AGEMA_signal_17203}), .b ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_17208, new_AGEMA_signal_17207, new_AGEMA_signal_17206}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_17439, new_AGEMA_signal_17438, new_AGEMA_signal_17437}), .b ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_17442, new_AGEMA_signal_17441, new_AGEMA_signal_17440}), .c ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_17445, new_AGEMA_signal_17444, new_AGEMA_signal_17443}), .b ({new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_17448, new_AGEMA_signal_17447, new_AGEMA_signal_17446}), .c ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_17217, new_AGEMA_signal_17216, new_AGEMA_signal_17215}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_17220, new_AGEMA_signal_17219, new_AGEMA_signal_17218}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_17217, new_AGEMA_signal_17216, new_AGEMA_signal_17215}), .b ({new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_17220, new_AGEMA_signal_17219, new_AGEMA_signal_17218}), .b ({new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_17451, new_AGEMA_signal_17450, new_AGEMA_signal_17449}), .b ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_17454, new_AGEMA_signal_17453, new_AGEMA_signal_17452}), .c ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_17457, new_AGEMA_signal_17456, new_AGEMA_signal_17455}), .b ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_17460, new_AGEMA_signal_17459, new_AGEMA_signal_17458}), .c ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_17229, new_AGEMA_signal_17228, new_AGEMA_signal_17227}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_17232, new_AGEMA_signal_17231, new_AGEMA_signal_17230}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_17229, new_AGEMA_signal_17228, new_AGEMA_signal_17227}), .b ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_17232, new_AGEMA_signal_17231, new_AGEMA_signal_17230}), .b ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_17463, new_AGEMA_signal_17462, new_AGEMA_signal_17461}), .b ({new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_17466, new_AGEMA_signal_17465, new_AGEMA_signal_17464}), .c ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_17469, new_AGEMA_signal_17468, new_AGEMA_signal_17467}), .b ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_17472, new_AGEMA_signal_17471, new_AGEMA_signal_17470}), .c ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_17241, new_AGEMA_signal_17240, new_AGEMA_signal_17239}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_17244, new_AGEMA_signal_17243, new_AGEMA_signal_17242}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_17241, new_AGEMA_signal_17240, new_AGEMA_signal_17239}), .b ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_17244, new_AGEMA_signal_17243, new_AGEMA_signal_17242}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_17475, new_AGEMA_signal_17474, new_AGEMA_signal_17473}), .b ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_17478, new_AGEMA_signal_17477, new_AGEMA_signal_17476}), .c ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_17481, new_AGEMA_signal_17480, new_AGEMA_signal_17479}), .b ({new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_17484, new_AGEMA_signal_17483, new_AGEMA_signal_17482}), .c ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_17253, new_AGEMA_signal_17252, new_AGEMA_signal_17251}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_17256, new_AGEMA_signal_17255, new_AGEMA_signal_17254}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_17253, new_AGEMA_signal_17252, new_AGEMA_signal_17251}), .b ({new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_17256, new_AGEMA_signal_17255, new_AGEMA_signal_17254}), .b ({new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_17487, new_AGEMA_signal_17486, new_AGEMA_signal_17485}), .b ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_17490, new_AGEMA_signal_17489, new_AGEMA_signal_17488}), .c ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_17493, new_AGEMA_signal_17492, new_AGEMA_signal_17491}), .b ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_17496, new_AGEMA_signal_17495, new_AGEMA_signal_17494}), .c ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_17265, new_AGEMA_signal_17264, new_AGEMA_signal_17263}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_17268, new_AGEMA_signal_17267, new_AGEMA_signal_17266}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_17265, new_AGEMA_signal_17264, new_AGEMA_signal_17263}), .b ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_17268, new_AGEMA_signal_17267, new_AGEMA_signal_17266}), .b ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_17499, new_AGEMA_signal_17498, new_AGEMA_signal_17497}), .b ({new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_17502, new_AGEMA_signal_17501, new_AGEMA_signal_17500}), .c ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_17505, new_AGEMA_signal_17504, new_AGEMA_signal_17503}), .b ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_17508, new_AGEMA_signal_17507, new_AGEMA_signal_17506}), .c ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_7562, new_AGEMA_signal_7561, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_17277, new_AGEMA_signal_17276, new_AGEMA_signal_17275}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_17280, new_AGEMA_signal_17279, new_AGEMA_signal_17278}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_17277, new_AGEMA_signal_17276, new_AGEMA_signal_17275}), .b ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_17280, new_AGEMA_signal_17279, new_AGEMA_signal_17278}), .b ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_17511, new_AGEMA_signal_17510, new_AGEMA_signal_17509}), .b ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_17514, new_AGEMA_signal_17513, new_AGEMA_signal_17512}), .c ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_17517, new_AGEMA_signal_17516, new_AGEMA_signal_17515}), .b ({new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_17520, new_AGEMA_signal_17519, new_AGEMA_signal_17518}), .c ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_17289, new_AGEMA_signal_17288, new_AGEMA_signal_17287}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_17292, new_AGEMA_signal_17291, new_AGEMA_signal_17290}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_17289, new_AGEMA_signal_17288, new_AGEMA_signal_17287}), .b ({new_AGEMA_signal_7574, new_AGEMA_signal_7573, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_17292, new_AGEMA_signal_17291, new_AGEMA_signal_17290}), .b ({new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_17523, new_AGEMA_signal_17522, new_AGEMA_signal_17521}), .b ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_17526, new_AGEMA_signal_17525, new_AGEMA_signal_17524}), .c ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_17529, new_AGEMA_signal_17528, new_AGEMA_signal_17527}), .b ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_17532, new_AGEMA_signal_17531, new_AGEMA_signal_17530}), .c ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_17301, new_AGEMA_signal_17300, new_AGEMA_signal_17299}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_7580, new_AGEMA_signal_7579, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_17304, new_AGEMA_signal_17303, new_AGEMA_signal_17302}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_17301, new_AGEMA_signal_17300, new_AGEMA_signal_17299}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_17304, new_AGEMA_signal_17303, new_AGEMA_signal_17302}), .b ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_17535, new_AGEMA_signal_17534, new_AGEMA_signal_17533}), .b ({new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_17538, new_AGEMA_signal_17537, new_AGEMA_signal_17536}), .c ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_17541, new_AGEMA_signal_17540, new_AGEMA_signal_17539}), .b ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_17544, new_AGEMA_signal_17543, new_AGEMA_signal_17542}), .c ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_7592, new_AGEMA_signal_7591, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_17313, new_AGEMA_signal_17312, new_AGEMA_signal_17311}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_17316, new_AGEMA_signal_17315, new_AGEMA_signal_17314}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_17313, new_AGEMA_signal_17312, new_AGEMA_signal_17311}), .b ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_17316, new_AGEMA_signal_17315, new_AGEMA_signal_17314}), .b ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_17547, new_AGEMA_signal_17546, new_AGEMA_signal_17545}), .b ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_17550, new_AGEMA_signal_17549, new_AGEMA_signal_17548}), .c ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_17553, new_AGEMA_signal_17552, new_AGEMA_signal_17551}), .b ({new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_17556, new_AGEMA_signal_17555, new_AGEMA_signal_17554}), .c ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_17325, new_AGEMA_signal_17324, new_AGEMA_signal_17323}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_17328, new_AGEMA_signal_17327, new_AGEMA_signal_17326}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_17325, new_AGEMA_signal_17324, new_AGEMA_signal_17323}), .b ({new_AGEMA_signal_7604, new_AGEMA_signal_7603, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_17328, new_AGEMA_signal_17327, new_AGEMA_signal_17326}), .b ({new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_17559, new_AGEMA_signal_17558, new_AGEMA_signal_17557}), .b ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_17562, new_AGEMA_signal_17561, new_AGEMA_signal_17560}), .c ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_17565, new_AGEMA_signal_17564, new_AGEMA_signal_17563}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_17568, new_AGEMA_signal_17567, new_AGEMA_signal_17566}), .c ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_17337, new_AGEMA_signal_17336, new_AGEMA_signal_17335}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_7610, new_AGEMA_signal_7609, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_17340, new_AGEMA_signal_17339, new_AGEMA_signal_17338}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_17337, new_AGEMA_signal_17336, new_AGEMA_signal_17335}), .b ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_17340, new_AGEMA_signal_17339, new_AGEMA_signal_17338}), .b ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_17571, new_AGEMA_signal_17570, new_AGEMA_signal_17569}), .b ({new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_17574, new_AGEMA_signal_17573, new_AGEMA_signal_17572}), .c ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_17577, new_AGEMA_signal_17576, new_AGEMA_signal_17575}), .b ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_17580, new_AGEMA_signal_17579, new_AGEMA_signal_17578}), .c ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_7622, new_AGEMA_signal_7621, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_17349, new_AGEMA_signal_17348, new_AGEMA_signal_17347}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_17352, new_AGEMA_signal_17351, new_AGEMA_signal_17350}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_17349, new_AGEMA_signal_17348, new_AGEMA_signal_17347}), .b ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_17352, new_AGEMA_signal_17351, new_AGEMA_signal_17350}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_17583, new_AGEMA_signal_17582, new_AGEMA_signal_17581}), .b ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_17586, new_AGEMA_signal_17585, new_AGEMA_signal_17584}), .c ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_17589, new_AGEMA_signal_17588, new_AGEMA_signal_17587}), .b ({new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_17592, new_AGEMA_signal_17591, new_AGEMA_signal_17590}), .c ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_17361, new_AGEMA_signal_17360, new_AGEMA_signal_17359}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_17364, new_AGEMA_signal_17363, new_AGEMA_signal_17362}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_17361, new_AGEMA_signal_17360, new_AGEMA_signal_17359}), .b ({new_AGEMA_signal_7634, new_AGEMA_signal_7633, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_17364, new_AGEMA_signal_17363, new_AGEMA_signal_17362}), .b ({new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_17595, new_AGEMA_signal_17594, new_AGEMA_signal_17593}), .b ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_17598, new_AGEMA_signal_17597, new_AGEMA_signal_17596}), .c ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_17601, new_AGEMA_signal_17600, new_AGEMA_signal_17599}), .b ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_17604, new_AGEMA_signal_17603, new_AGEMA_signal_17602}), .c ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_7442, new_AGEMA_signal_7441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_17373, new_AGEMA_signal_17372, new_AGEMA_signal_17371}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_17376, new_AGEMA_signal_17375, new_AGEMA_signal_17374}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_17373, new_AGEMA_signal_17372, new_AGEMA_signal_17371}), .b ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_17376, new_AGEMA_signal_17375, new_AGEMA_signal_17374}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_17607, new_AGEMA_signal_17606, new_AGEMA_signal_17605}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_17610, new_AGEMA_signal_17609, new_AGEMA_signal_17608}), .c ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_17613, new_AGEMA_signal_17612, new_AGEMA_signal_17611}), .b ({new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_17616, new_AGEMA_signal_17615, new_AGEMA_signal_17614}), .c ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_17385, new_AGEMA_signal_17384, new_AGEMA_signal_17383}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_17388, new_AGEMA_signal_17387, new_AGEMA_signal_17386}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_17385, new_AGEMA_signal_17384, new_AGEMA_signal_17383}), .b ({new_AGEMA_signal_7454, new_AGEMA_signal_7453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_17388, new_AGEMA_signal_17387, new_AGEMA_signal_17386}), .b ({new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_17619, new_AGEMA_signal_17618, new_AGEMA_signal_17617}), .b ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_17622, new_AGEMA_signal_17621, new_AGEMA_signal_17620}), .c ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_17625, new_AGEMA_signal_17624, new_AGEMA_signal_17623}), .b ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_17628, new_AGEMA_signal_17627, new_AGEMA_signal_17626}), .c ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_17397, new_AGEMA_signal_17396, new_AGEMA_signal_17395}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_7460, new_AGEMA_signal_7459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_17400, new_AGEMA_signal_17399, new_AGEMA_signal_17398}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_17397, new_AGEMA_signal_17396, new_AGEMA_signal_17395}), .b ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_17400, new_AGEMA_signal_17399, new_AGEMA_signal_17398}), .b ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_17631, new_AGEMA_signal_17630, new_AGEMA_signal_17629}), .b ({new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_17634, new_AGEMA_signal_17633, new_AGEMA_signal_17632}), .c ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_17637, new_AGEMA_signal_17636, new_AGEMA_signal_17635}), .b ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_17640, new_AGEMA_signal_17639, new_AGEMA_signal_17638}), .c ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_7472, new_AGEMA_signal_7471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_17409, new_AGEMA_signal_17408, new_AGEMA_signal_17407}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_17412, new_AGEMA_signal_17411, new_AGEMA_signal_17410}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_7670, new_AGEMA_signal_7669, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_17409, new_AGEMA_signal_17408, new_AGEMA_signal_17407}), .b ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_17412, new_AGEMA_signal_17411, new_AGEMA_signal_17410}), .b ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_17643, new_AGEMA_signal_17642, new_AGEMA_signal_17641}), .b ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_17646, new_AGEMA_signal_17645, new_AGEMA_signal_17644}), .c ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_17649, new_AGEMA_signal_17648, new_AGEMA_signal_17647}), .b ({new_AGEMA_signal_7670, new_AGEMA_signal_7669, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_17652, new_AGEMA_signal_17651, new_AGEMA_signal_17650}), .c ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (new_AGEMA_signal_17173), .Q (new_AGEMA_signal_17413) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_17174), .Q (new_AGEMA_signal_17414) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_17175), .Q (new_AGEMA_signal_17415) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_17416) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_7485), .Q (new_AGEMA_signal_17417) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_17418) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_17176), .Q (new_AGEMA_signal_17419) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_17177), .Q (new_AGEMA_signal_17420) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (new_AGEMA_signal_17178), .Q (new_AGEMA_signal_17421) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_17422) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_7685), .Q (new_AGEMA_signal_17423) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_7686), .Q (new_AGEMA_signal_17424) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (new_AGEMA_signal_17185), .Q (new_AGEMA_signal_17425) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_17186), .Q (new_AGEMA_signal_17426) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_17187), .Q (new_AGEMA_signal_17427) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_17428) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_17429) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_17430) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_17188), .Q (new_AGEMA_signal_17431) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_17189), .Q (new_AGEMA_signal_17432) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_17190), .Q (new_AGEMA_signal_17433) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_17434) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_7695), .Q (new_AGEMA_signal_17435) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_17436) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (new_AGEMA_signal_17197), .Q (new_AGEMA_signal_17437) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_17198), .Q (new_AGEMA_signal_17438) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_17199), .Q (new_AGEMA_signal_17439) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_17440) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_7505), .Q (new_AGEMA_signal_17441) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_7506), .Q (new_AGEMA_signal_17442) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_17200), .Q (new_AGEMA_signal_17443) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_17201), .Q (new_AGEMA_signal_17444) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (new_AGEMA_signal_17202), .Q (new_AGEMA_signal_17445) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_17446) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_7705), .Q (new_AGEMA_signal_17447) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_7706), .Q (new_AGEMA_signal_17448) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (new_AGEMA_signal_17209), .Q (new_AGEMA_signal_17449) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_17210), .Q (new_AGEMA_signal_17450) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_17211), .Q (new_AGEMA_signal_17451) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_17452) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_17453) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_17454) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_17212), .Q (new_AGEMA_signal_17455) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_17213), .Q (new_AGEMA_signal_17456) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_17214), .Q (new_AGEMA_signal_17457) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_17458) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_7715), .Q (new_AGEMA_signal_17459) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_7716), .Q (new_AGEMA_signal_17460) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (new_AGEMA_signal_17221), .Q (new_AGEMA_signal_17461) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_17222), .Q (new_AGEMA_signal_17462) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_17223), .Q (new_AGEMA_signal_17463) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M33), .Q (new_AGEMA_signal_17464) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_7525), .Q (new_AGEMA_signal_17465) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_17466) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_17224), .Q (new_AGEMA_signal_17467) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_17225), .Q (new_AGEMA_signal_17468) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (new_AGEMA_signal_17226), .Q (new_AGEMA_signal_17469) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (SubBytesIns_Inst_Sbox_4_M36), .Q (new_AGEMA_signal_17470) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_7725), .Q (new_AGEMA_signal_17471) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_7726), .Q (new_AGEMA_signal_17472) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (new_AGEMA_signal_17233), .Q (new_AGEMA_signal_17473) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_17234), .Q (new_AGEMA_signal_17474) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_17235), .Q (new_AGEMA_signal_17475) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M33), .Q (new_AGEMA_signal_17476) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_17477) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_17478) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_17236), .Q (new_AGEMA_signal_17479) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_17237), .Q (new_AGEMA_signal_17480) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (new_AGEMA_signal_17238), .Q (new_AGEMA_signal_17481) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (SubBytesIns_Inst_Sbox_5_M36), .Q (new_AGEMA_signal_17482) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_17483) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_17484) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C (clk), .D (new_AGEMA_signal_17245), .Q (new_AGEMA_signal_17485) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_17246), .Q (new_AGEMA_signal_17486) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_17247), .Q (new_AGEMA_signal_17487) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M33), .Q (new_AGEMA_signal_17488) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C (clk), .D (new_AGEMA_signal_7545), .Q (new_AGEMA_signal_17489) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_7546), .Q (new_AGEMA_signal_17490) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_17248), .Q (new_AGEMA_signal_17491) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_17249), .Q (new_AGEMA_signal_17492) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C (clk), .D (new_AGEMA_signal_17250), .Q (new_AGEMA_signal_17493) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C (clk), .D (SubBytesIns_Inst_Sbox_6_M36), .Q (new_AGEMA_signal_17494) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_7745), .Q (new_AGEMA_signal_17495) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_7746), .Q (new_AGEMA_signal_17496) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C (clk), .D (new_AGEMA_signal_17257), .Q (new_AGEMA_signal_17497) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_17258), .Q (new_AGEMA_signal_17498) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_17259), .Q (new_AGEMA_signal_17499) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M33), .Q (new_AGEMA_signal_17500) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C (clk), .D (new_AGEMA_signal_7555), .Q (new_AGEMA_signal_17501) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_17502) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_17260), .Q (new_AGEMA_signal_17503) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_17261), .Q (new_AGEMA_signal_17504) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C (clk), .D (new_AGEMA_signal_17262), .Q (new_AGEMA_signal_17505) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C (clk), .D (SubBytesIns_Inst_Sbox_7_M36), .Q (new_AGEMA_signal_17506) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_7755), .Q (new_AGEMA_signal_17507) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_17508) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C (clk), .D (new_AGEMA_signal_17269), .Q (new_AGEMA_signal_17509) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_17270), .Q (new_AGEMA_signal_17510) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_17271), .Q (new_AGEMA_signal_17511) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M33), .Q (new_AGEMA_signal_17512) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C (clk), .D (new_AGEMA_signal_7565), .Q (new_AGEMA_signal_17513) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_7566), .Q (new_AGEMA_signal_17514) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_17272), .Q (new_AGEMA_signal_17515) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_17273), .Q (new_AGEMA_signal_17516) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C (clk), .D (new_AGEMA_signal_17274), .Q (new_AGEMA_signal_17517) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C (clk), .D (SubBytesIns_Inst_Sbox_8_M36), .Q (new_AGEMA_signal_17518) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_7765), .Q (new_AGEMA_signal_17519) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_7766), .Q (new_AGEMA_signal_17520) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C (clk), .D (new_AGEMA_signal_17281), .Q (new_AGEMA_signal_17521) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_17282), .Q (new_AGEMA_signal_17522) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_17283), .Q (new_AGEMA_signal_17523) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M33), .Q (new_AGEMA_signal_17524) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_17525) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_17526) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_17284), .Q (new_AGEMA_signal_17527) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_17285), .Q (new_AGEMA_signal_17528) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C (clk), .D (new_AGEMA_signal_17286), .Q (new_AGEMA_signal_17529) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C (clk), .D (SubBytesIns_Inst_Sbox_9_M36), .Q (new_AGEMA_signal_17530) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_17531) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_7776), .Q (new_AGEMA_signal_17532) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C (clk), .D (new_AGEMA_signal_17293), .Q (new_AGEMA_signal_17533) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_17294), .Q (new_AGEMA_signal_17534) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_17295), .Q (new_AGEMA_signal_17535) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M33), .Q (new_AGEMA_signal_17536) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C (clk), .D (new_AGEMA_signal_7585), .Q (new_AGEMA_signal_17537) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_7586), .Q (new_AGEMA_signal_17538) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_17296), .Q (new_AGEMA_signal_17539) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_17297), .Q (new_AGEMA_signal_17540) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C (clk), .D (new_AGEMA_signal_17298), .Q (new_AGEMA_signal_17541) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C (clk), .D (SubBytesIns_Inst_Sbox_10_M36), .Q (new_AGEMA_signal_17542) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_7785), .Q (new_AGEMA_signal_17543) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_7786), .Q (new_AGEMA_signal_17544) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C (clk), .D (new_AGEMA_signal_17305), .Q (new_AGEMA_signal_17545) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_17306), .Q (new_AGEMA_signal_17546) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_17307), .Q (new_AGEMA_signal_17547) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M33), .Q (new_AGEMA_signal_17548) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C (clk), .D (new_AGEMA_signal_7595), .Q (new_AGEMA_signal_17549) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_17550) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_17308), .Q (new_AGEMA_signal_17551) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_17309), .Q (new_AGEMA_signal_17552) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C (clk), .D (new_AGEMA_signal_17310), .Q (new_AGEMA_signal_17553) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C (clk), .D (SubBytesIns_Inst_Sbox_11_M36), .Q (new_AGEMA_signal_17554) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_7795), .Q (new_AGEMA_signal_17555) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_17556) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C (clk), .D (new_AGEMA_signal_17317), .Q (new_AGEMA_signal_17557) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_17318), .Q (new_AGEMA_signal_17558) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_17319), .Q (new_AGEMA_signal_17559) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M33), .Q (new_AGEMA_signal_17560) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C (clk), .D (new_AGEMA_signal_7605), .Q (new_AGEMA_signal_17561) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_7606), .Q (new_AGEMA_signal_17562) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_17320), .Q (new_AGEMA_signal_17563) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_17321), .Q (new_AGEMA_signal_17564) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C (clk), .D (new_AGEMA_signal_17322), .Q (new_AGEMA_signal_17565) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C (clk), .D (SubBytesIns_Inst_Sbox_12_M36), .Q (new_AGEMA_signal_17566) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_17567) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_7806), .Q (new_AGEMA_signal_17568) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C (clk), .D (new_AGEMA_signal_17329), .Q (new_AGEMA_signal_17569) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_17330), .Q (new_AGEMA_signal_17570) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_17331), .Q (new_AGEMA_signal_17571) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M33), .Q (new_AGEMA_signal_17572) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_17573) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_17574) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_17332), .Q (new_AGEMA_signal_17575) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_17333), .Q (new_AGEMA_signal_17576) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C (clk), .D (new_AGEMA_signal_17334), .Q (new_AGEMA_signal_17577) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C (clk), .D (SubBytesIns_Inst_Sbox_13_M36), .Q (new_AGEMA_signal_17578) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_7815), .Q (new_AGEMA_signal_17579) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_17580) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C (clk), .D (new_AGEMA_signal_17341), .Q (new_AGEMA_signal_17581) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_17342), .Q (new_AGEMA_signal_17582) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_17343), .Q (new_AGEMA_signal_17583) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M33), .Q (new_AGEMA_signal_17584) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C (clk), .D (new_AGEMA_signal_7625), .Q (new_AGEMA_signal_17585) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_7626), .Q (new_AGEMA_signal_17586) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_17344), .Q (new_AGEMA_signal_17587) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_17345), .Q (new_AGEMA_signal_17588) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C (clk), .D (new_AGEMA_signal_17346), .Q (new_AGEMA_signal_17589) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C (clk), .D (SubBytesIns_Inst_Sbox_14_M36), .Q (new_AGEMA_signal_17590) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_7825), .Q (new_AGEMA_signal_17591) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_7826), .Q (new_AGEMA_signal_17592) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C (clk), .D (new_AGEMA_signal_17353), .Q (new_AGEMA_signal_17593) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_17354), .Q (new_AGEMA_signal_17594) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_17355), .Q (new_AGEMA_signal_17595) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M33), .Q (new_AGEMA_signal_17596) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C (clk), .D (new_AGEMA_signal_7635), .Q (new_AGEMA_signal_17597) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_17598) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_17356), .Q (new_AGEMA_signal_17599) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_17357), .Q (new_AGEMA_signal_17600) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C (clk), .D (new_AGEMA_signal_17358), .Q (new_AGEMA_signal_17601) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C (clk), .D (SubBytesIns_Inst_Sbox_15_M36), .Q (new_AGEMA_signal_17602) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_17603) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_17604) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C (clk), .D (new_AGEMA_signal_17365), .Q (new_AGEMA_signal_17605) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_17366), .Q (new_AGEMA_signal_17606) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_17367), .Q (new_AGEMA_signal_17607) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_17608) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C (clk), .D (new_AGEMA_signal_7445), .Q (new_AGEMA_signal_17609) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_17610) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_17368), .Q (new_AGEMA_signal_17611) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_17369), .Q (new_AGEMA_signal_17612) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C (clk), .D (new_AGEMA_signal_17370), .Q (new_AGEMA_signal_17613) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_17614) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_17615) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_7646), .Q (new_AGEMA_signal_17616) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C (clk), .D (new_AGEMA_signal_17377), .Q (new_AGEMA_signal_17617) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_17378), .Q (new_AGEMA_signal_17618) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_17379), .Q (new_AGEMA_signal_17619) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_17620) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_17621) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_17622) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_17380), .Q (new_AGEMA_signal_17623) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_17381), .Q (new_AGEMA_signal_17624) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C (clk), .D (new_AGEMA_signal_17382), .Q (new_AGEMA_signal_17625) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_17626) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_17627) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_7656), .Q (new_AGEMA_signal_17628) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C (clk), .D (new_AGEMA_signal_17389), .Q (new_AGEMA_signal_17629) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_17390), .Q (new_AGEMA_signal_17630) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_17391), .Q (new_AGEMA_signal_17631) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_17632) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C (clk), .D (new_AGEMA_signal_7465), .Q (new_AGEMA_signal_17633) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_7466), .Q (new_AGEMA_signal_17634) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_17392), .Q (new_AGEMA_signal_17635) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_17393), .Q (new_AGEMA_signal_17636) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C (clk), .D (new_AGEMA_signal_17394), .Q (new_AGEMA_signal_17637) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_17638) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_7665), .Q (new_AGEMA_signal_17639) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_7666), .Q (new_AGEMA_signal_17640) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C (clk), .D (new_AGEMA_signal_17401), .Q (new_AGEMA_signal_17641) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_17402), .Q (new_AGEMA_signal_17642) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_17403), .Q (new_AGEMA_signal_17643) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_17644) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_17645) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_17646) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_17404), .Q (new_AGEMA_signal_17647) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_17405), .Q (new_AGEMA_signal_17648) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C (clk), .D (new_AGEMA_signal_17406), .Q (new_AGEMA_signal_17649) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C (clk), .D (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_17650) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_7675), .Q (new_AGEMA_signal_17651) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_17652) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_17654), .Q (new_AGEMA_signal_17655) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_17658), .Q (new_AGEMA_signal_17659) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_17662), .Q (new_AGEMA_signal_17663) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_17666), .Q (new_AGEMA_signal_17667) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_17670), .Q (new_AGEMA_signal_17671) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_17674), .Q (new_AGEMA_signal_17675) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_17678), .Q (new_AGEMA_signal_17679) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_17682), .Q (new_AGEMA_signal_17683) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_17686), .Q (new_AGEMA_signal_17687) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_17690), .Q (new_AGEMA_signal_17691) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_17694), .Q (new_AGEMA_signal_17695) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_17698), .Q (new_AGEMA_signal_17699) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_17702), .Q (new_AGEMA_signal_17703) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_17706), .Q (new_AGEMA_signal_17707) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_17710), .Q (new_AGEMA_signal_17711) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_17714), .Q (new_AGEMA_signal_17715) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_17718), .Q (new_AGEMA_signal_17719) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_17722), .Q (new_AGEMA_signal_17723) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_17726), .Q (new_AGEMA_signal_17727) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_17730), .Q (new_AGEMA_signal_17731) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_17734), .Q (new_AGEMA_signal_17735) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_17738), .Q (new_AGEMA_signal_17739) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_17742), .Q (new_AGEMA_signal_17743) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_17746), .Q (new_AGEMA_signal_17747) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_17750), .Q (new_AGEMA_signal_17751) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_17754), .Q (new_AGEMA_signal_17755) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_17758), .Q (new_AGEMA_signal_17759) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_17762), .Q (new_AGEMA_signal_17763) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_17766), .Q (new_AGEMA_signal_17767) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_17770), .Q (new_AGEMA_signal_17771) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_17774), .Q (new_AGEMA_signal_17775) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_17778), .Q (new_AGEMA_signal_17779) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_17782), .Q (new_AGEMA_signal_17783) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_17786), .Q (new_AGEMA_signal_17787) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_17790), .Q (new_AGEMA_signal_17791) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_17794), .Q (new_AGEMA_signal_17795) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_17798), .Q (new_AGEMA_signal_17799) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_17802), .Q (new_AGEMA_signal_17803) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_17806), .Q (new_AGEMA_signal_17807) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_17810), .Q (new_AGEMA_signal_17811) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_17814), .Q (new_AGEMA_signal_17815) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_17818), .Q (new_AGEMA_signal_17819) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_17822), .Q (new_AGEMA_signal_17823) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_17826), .Q (new_AGEMA_signal_17827) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_17830), .Q (new_AGEMA_signal_17831) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_17834), .Q (new_AGEMA_signal_17835) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_17838), .Q (new_AGEMA_signal_17839) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_17842), .Q (new_AGEMA_signal_17843) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_17846), .Q (new_AGEMA_signal_17847) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_17850), .Q (new_AGEMA_signal_17851) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_17854), .Q (new_AGEMA_signal_17855) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_17858), .Q (new_AGEMA_signal_17859) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_17862), .Q (new_AGEMA_signal_17863) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_17866), .Q (new_AGEMA_signal_17867) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_17870), .Q (new_AGEMA_signal_17871) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_17874), .Q (new_AGEMA_signal_17875) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_17878), .Q (new_AGEMA_signal_17879) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_17882), .Q (new_AGEMA_signal_17883) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_17886), .Q (new_AGEMA_signal_17887) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_17890), .Q (new_AGEMA_signal_17891) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_17894), .Q (new_AGEMA_signal_17895) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_17898), .Q (new_AGEMA_signal_17899) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_17902), .Q (new_AGEMA_signal_17903) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_17906), .Q (new_AGEMA_signal_17907) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_17910), .Q (new_AGEMA_signal_17911) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_17914), .Q (new_AGEMA_signal_17915) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_17918), .Q (new_AGEMA_signal_17919) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_17922), .Q (new_AGEMA_signal_17923) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_17926), .Q (new_AGEMA_signal_17927) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_17930), .Q (new_AGEMA_signal_17931) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_17934), .Q (new_AGEMA_signal_17935) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_17938), .Q (new_AGEMA_signal_17939) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_17942), .Q (new_AGEMA_signal_17943) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_17946), .Q (new_AGEMA_signal_17947) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_17950), .Q (new_AGEMA_signal_17951) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_17954), .Q (new_AGEMA_signal_17955) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_17958), .Q (new_AGEMA_signal_17959) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_17962), .Q (new_AGEMA_signal_17963) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_17966), .Q (new_AGEMA_signal_17967) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_17970), .Q (new_AGEMA_signal_17971) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_17974), .Q (new_AGEMA_signal_17975) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_17978), .Q (new_AGEMA_signal_17979) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_17982), .Q (new_AGEMA_signal_17983) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_17986), .Q (new_AGEMA_signal_17987) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_17990), .Q (new_AGEMA_signal_17991) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_17994), .Q (new_AGEMA_signal_17995) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_17998), .Q (new_AGEMA_signal_17999) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_18002), .Q (new_AGEMA_signal_18003) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_18006), .Q (new_AGEMA_signal_18007) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_18010), .Q (new_AGEMA_signal_18011) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_18014), .Q (new_AGEMA_signal_18015) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_18018), .Q (new_AGEMA_signal_18019) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_18022), .Q (new_AGEMA_signal_18023) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_18026), .Q (new_AGEMA_signal_18027) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_18030), .Q (new_AGEMA_signal_18031) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_18034), .Q (new_AGEMA_signal_18035) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_18038), .Q (new_AGEMA_signal_18039) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_18042), .Q (new_AGEMA_signal_18043) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_18046), .Q (new_AGEMA_signal_18047) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_18050), .Q (new_AGEMA_signal_18051) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_18054), .Q (new_AGEMA_signal_18055) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_18058), .Q (new_AGEMA_signal_18059) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_18062), .Q (new_AGEMA_signal_18063) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_18066), .Q (new_AGEMA_signal_18067) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_18070), .Q (new_AGEMA_signal_18071) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_18074), .Q (new_AGEMA_signal_18075) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_18078), .Q (new_AGEMA_signal_18079) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_18082), .Q (new_AGEMA_signal_18083) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_18086), .Q (new_AGEMA_signal_18087) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_18090), .Q (new_AGEMA_signal_18091) ) ;
    buf_clk new_AGEMA_reg_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_18094), .Q (new_AGEMA_signal_18095) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_18098), .Q (new_AGEMA_signal_18099) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_18102), .Q (new_AGEMA_signal_18103) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_18106), .Q (new_AGEMA_signal_18107) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_18110), .Q (new_AGEMA_signal_18111) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_18114), .Q (new_AGEMA_signal_18115) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_18118), .Q (new_AGEMA_signal_18119) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_18122), .Q (new_AGEMA_signal_18123) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_18126), .Q (new_AGEMA_signal_18127) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_18130), .Q (new_AGEMA_signal_18131) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_18134), .Q (new_AGEMA_signal_18135) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_18138), .Q (new_AGEMA_signal_18139) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_18142), .Q (new_AGEMA_signal_18143) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_18146), .Q (new_AGEMA_signal_18147) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_18150), .Q (new_AGEMA_signal_18151) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_18154), .Q (new_AGEMA_signal_18155) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_18158), .Q (new_AGEMA_signal_18159) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_18162), .Q (new_AGEMA_signal_18163) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_18166), .Q (new_AGEMA_signal_18167) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_18170), .Q (new_AGEMA_signal_18171) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_18174), .Q (new_AGEMA_signal_18175) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_18178), .Q (new_AGEMA_signal_18179) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_18182), .Q (new_AGEMA_signal_18183) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_18186), .Q (new_AGEMA_signal_18187) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_18190), .Q (new_AGEMA_signal_18191) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_18194), .Q (new_AGEMA_signal_18195) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_18198), .Q (new_AGEMA_signal_18199) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_18202), .Q (new_AGEMA_signal_18203) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_18206), .Q (new_AGEMA_signal_18207) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_18210), .Q (new_AGEMA_signal_18211) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_18214), .Q (new_AGEMA_signal_18215) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_18218), .Q (new_AGEMA_signal_18219) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_18222), .Q (new_AGEMA_signal_18223) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_18226), .Q (new_AGEMA_signal_18227) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_18230), .Q (new_AGEMA_signal_18231) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_18234), .Q (new_AGEMA_signal_18235) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_18238), .Q (new_AGEMA_signal_18239) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_18242), .Q (new_AGEMA_signal_18243) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_18246), .Q (new_AGEMA_signal_18247) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_18250), .Q (new_AGEMA_signal_18251) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_18254), .Q (new_AGEMA_signal_18255) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_18258), .Q (new_AGEMA_signal_18259) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_18262), .Q (new_AGEMA_signal_18263) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_18266), .Q (new_AGEMA_signal_18267) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_18270), .Q (new_AGEMA_signal_18271) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_18274), .Q (new_AGEMA_signal_18275) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_18278), .Q (new_AGEMA_signal_18279) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_18282), .Q (new_AGEMA_signal_18283) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_18286), .Q (new_AGEMA_signal_18287) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_18290), .Q (new_AGEMA_signal_18291) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_18294), .Q (new_AGEMA_signal_18295) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_18298), .Q (new_AGEMA_signal_18299) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_18302), .Q (new_AGEMA_signal_18303) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_18306), .Q (new_AGEMA_signal_18307) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_18310), .Q (new_AGEMA_signal_18311) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_18314), .Q (new_AGEMA_signal_18315) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_18318), .Q (new_AGEMA_signal_18319) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_18322), .Q (new_AGEMA_signal_18323) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_18326), .Q (new_AGEMA_signal_18327) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_18330), .Q (new_AGEMA_signal_18331) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_18334), .Q (new_AGEMA_signal_18335) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_18338), .Q (new_AGEMA_signal_18339) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_18342), .Q (new_AGEMA_signal_18343) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_18346), .Q (new_AGEMA_signal_18347) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_18350), .Q (new_AGEMA_signal_18351) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_18354), .Q (new_AGEMA_signal_18355) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_18358), .Q (new_AGEMA_signal_18359) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_18362), .Q (new_AGEMA_signal_18363) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_18366), .Q (new_AGEMA_signal_18367) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_18370), .Q (new_AGEMA_signal_18371) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_18374), .Q (new_AGEMA_signal_18375) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_18378), .Q (new_AGEMA_signal_18379) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_18382), .Q (new_AGEMA_signal_18383) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_18386), .Q (new_AGEMA_signal_18387) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_18390), .Q (new_AGEMA_signal_18391) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_18394), .Q (new_AGEMA_signal_18395) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_18398), .Q (new_AGEMA_signal_18399) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_18402), .Q (new_AGEMA_signal_18403) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_18406), .Q (new_AGEMA_signal_18407) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_18410), .Q (new_AGEMA_signal_18411) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_18414), .Q (new_AGEMA_signal_18415) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_18418), .Q (new_AGEMA_signal_18419) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_18422), .Q (new_AGEMA_signal_18423) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_18426), .Q (new_AGEMA_signal_18427) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_18430), .Q (new_AGEMA_signal_18431) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_18434), .Q (new_AGEMA_signal_18435) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_18438), .Q (new_AGEMA_signal_18439) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_18442), .Q (new_AGEMA_signal_18443) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_18446), .Q (new_AGEMA_signal_18447) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_18450), .Q (new_AGEMA_signal_18451) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_18454), .Q (new_AGEMA_signal_18455) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_18458), .Q (new_AGEMA_signal_18459) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_18462), .Q (new_AGEMA_signal_18463) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_18466), .Q (new_AGEMA_signal_18467) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_18470), .Q (new_AGEMA_signal_18471) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_18474), .Q (new_AGEMA_signal_18475) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_18478), .Q (new_AGEMA_signal_18479) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_18482), .Q (new_AGEMA_signal_18483) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_18486), .Q (new_AGEMA_signal_18487) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_18490), .Q (new_AGEMA_signal_18491) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_18494), .Q (new_AGEMA_signal_18495) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_18498), .Q (new_AGEMA_signal_18499) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_18502), .Q (new_AGEMA_signal_18503) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_18506), .Q (new_AGEMA_signal_18507) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_18510), .Q (new_AGEMA_signal_18511) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_18514), .Q (new_AGEMA_signal_18515) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_18518), .Q (new_AGEMA_signal_18519) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_18522), .Q (new_AGEMA_signal_18523) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_18526), .Q (new_AGEMA_signal_18527) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_18530), .Q (new_AGEMA_signal_18531) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_18534), .Q (new_AGEMA_signal_18535) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_18538), .Q (new_AGEMA_signal_18539) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_18542), .Q (new_AGEMA_signal_18543) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_18546), .Q (new_AGEMA_signal_18547) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_18550), .Q (new_AGEMA_signal_18551) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_18554), .Q (new_AGEMA_signal_18555) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_18558), .Q (new_AGEMA_signal_18559) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_18562), .Q (new_AGEMA_signal_18563) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_18566), .Q (new_AGEMA_signal_18567) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_18570), .Q (new_AGEMA_signal_18571) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_18574), .Q (new_AGEMA_signal_18575) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_18578), .Q (new_AGEMA_signal_18579) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_18582), .Q (new_AGEMA_signal_18583) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_18586), .Q (new_AGEMA_signal_18587) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_18590), .Q (new_AGEMA_signal_18591) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_18594), .Q (new_AGEMA_signal_18595) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_18598), .Q (new_AGEMA_signal_18599) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_18602), .Q (new_AGEMA_signal_18603) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_18606), .Q (new_AGEMA_signal_18607) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_18610), .Q (new_AGEMA_signal_18611) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_18614), .Q (new_AGEMA_signal_18615) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_18618), .Q (new_AGEMA_signal_18619) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_18622), .Q (new_AGEMA_signal_18623) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_18626), .Q (new_AGEMA_signal_18627) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_18630), .Q (new_AGEMA_signal_18631) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_18634), .Q (new_AGEMA_signal_18635) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_18638), .Q (new_AGEMA_signal_18639) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_18642), .Q (new_AGEMA_signal_18643) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_18646), .Q (new_AGEMA_signal_18647) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_18650), .Q (new_AGEMA_signal_18651) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_18654), .Q (new_AGEMA_signal_18655) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_18658), .Q (new_AGEMA_signal_18659) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_18662), .Q (new_AGEMA_signal_18663) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_18666), .Q (new_AGEMA_signal_18667) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_18670), .Q (new_AGEMA_signal_18671) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_18674), .Q (new_AGEMA_signal_18675) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_18678), .Q (new_AGEMA_signal_18679) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_18682), .Q (new_AGEMA_signal_18683) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_18686), .Q (new_AGEMA_signal_18687) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_18690), .Q (new_AGEMA_signal_18691) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_18694), .Q (new_AGEMA_signal_18695) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_18698), .Q (new_AGEMA_signal_18699) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_18702), .Q (new_AGEMA_signal_18703) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_18706), .Q (new_AGEMA_signal_18707) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_18710), .Q (new_AGEMA_signal_18711) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_18714), .Q (new_AGEMA_signal_18715) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_18718), .Q (new_AGEMA_signal_18719) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_18722), .Q (new_AGEMA_signal_18723) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_18726), .Q (new_AGEMA_signal_18727) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_18730), .Q (new_AGEMA_signal_18731) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_18734), .Q (new_AGEMA_signal_18735) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_18738), .Q (new_AGEMA_signal_18739) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_18742), .Q (new_AGEMA_signal_18743) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_18746), .Q (new_AGEMA_signal_18747) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_18750), .Q (new_AGEMA_signal_18751) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_18754), .Q (new_AGEMA_signal_18755) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_18758), .Q (new_AGEMA_signal_18759) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_18762), .Q (new_AGEMA_signal_18763) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_18766), .Q (new_AGEMA_signal_18767) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_18770), .Q (new_AGEMA_signal_18771) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C (clk), .D (new_AGEMA_signal_18774), .Q (new_AGEMA_signal_18775) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_18778), .Q (new_AGEMA_signal_18779) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_18782), .Q (new_AGEMA_signal_18783) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C (clk), .D (new_AGEMA_signal_18786), .Q (new_AGEMA_signal_18787) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_18790), .Q (new_AGEMA_signal_18791) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_18794), .Q (new_AGEMA_signal_18795) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C (clk), .D (new_AGEMA_signal_18798), .Q (new_AGEMA_signal_18799) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_18802), .Q (new_AGEMA_signal_18803) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_18806), .Q (new_AGEMA_signal_18807) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C (clk), .D (new_AGEMA_signal_18810), .Q (new_AGEMA_signal_18811) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_18814), .Q (new_AGEMA_signal_18815) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_18818), .Q (new_AGEMA_signal_18819) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C (clk), .D (new_AGEMA_signal_18822), .Q (new_AGEMA_signal_18823) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_18826), .Q (new_AGEMA_signal_18827) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_18830), .Q (new_AGEMA_signal_18831) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C (clk), .D (new_AGEMA_signal_18834), .Q (new_AGEMA_signal_18835) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_18838), .Q (new_AGEMA_signal_18839) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_18842), .Q (new_AGEMA_signal_18843) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C (clk), .D (new_AGEMA_signal_18846), .Q (new_AGEMA_signal_18847) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_18850), .Q (new_AGEMA_signal_18851) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_18854), .Q (new_AGEMA_signal_18855) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C (clk), .D (new_AGEMA_signal_18858), .Q (new_AGEMA_signal_18859) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_18862), .Q (new_AGEMA_signal_18863) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_18866), .Q (new_AGEMA_signal_18867) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C (clk), .D (new_AGEMA_signal_18870), .Q (new_AGEMA_signal_18871) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_18874), .Q (new_AGEMA_signal_18875) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_18878), .Q (new_AGEMA_signal_18879) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C (clk), .D (new_AGEMA_signal_18882), .Q (new_AGEMA_signal_18883) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_18886), .Q (new_AGEMA_signal_18887) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_18890), .Q (new_AGEMA_signal_18891) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C (clk), .D (new_AGEMA_signal_18894), .Q (new_AGEMA_signal_18895) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_18898), .Q (new_AGEMA_signal_18899) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C (clk), .D (new_AGEMA_signal_18902), .Q (new_AGEMA_signal_18903) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C (clk), .D (new_AGEMA_signal_18906), .Q (new_AGEMA_signal_18907) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_18910), .Q (new_AGEMA_signal_18911) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_18914), .Q (new_AGEMA_signal_18915) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C (clk), .D (new_AGEMA_signal_18918), .Q (new_AGEMA_signal_18919) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_18922), .Q (new_AGEMA_signal_18923) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_18926), .Q (new_AGEMA_signal_18927) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C (clk), .D (new_AGEMA_signal_18930), .Q (new_AGEMA_signal_18931) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_18934), .Q (new_AGEMA_signal_18935) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C (clk), .D (new_AGEMA_signal_18938), .Q (new_AGEMA_signal_18939) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C (clk), .D (new_AGEMA_signal_18942), .Q (new_AGEMA_signal_18943) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_18946), .Q (new_AGEMA_signal_18947) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_18950), .Q (new_AGEMA_signal_18951) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C (clk), .D (new_AGEMA_signal_18954), .Q (new_AGEMA_signal_18955) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_18958), .Q (new_AGEMA_signal_18959) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_18962), .Q (new_AGEMA_signal_18963) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C (clk), .D (new_AGEMA_signal_18966), .Q (new_AGEMA_signal_18967) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_18970), .Q (new_AGEMA_signal_18971) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C (clk), .D (new_AGEMA_signal_18974), .Q (new_AGEMA_signal_18975) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C (clk), .D (new_AGEMA_signal_18978), .Q (new_AGEMA_signal_18979) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_18982), .Q (new_AGEMA_signal_18983) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_18986), .Q (new_AGEMA_signal_18987) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C (clk), .D (new_AGEMA_signal_18990), .Q (new_AGEMA_signal_18991) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_18994), .Q (new_AGEMA_signal_18995) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_18998), .Q (new_AGEMA_signal_18999) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C (clk), .D (new_AGEMA_signal_19002), .Q (new_AGEMA_signal_19003) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_19006), .Q (new_AGEMA_signal_19007) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C (clk), .D (new_AGEMA_signal_19010), .Q (new_AGEMA_signal_19011) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C (clk), .D (new_AGEMA_signal_19014), .Q (new_AGEMA_signal_19015) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_19018), .Q (new_AGEMA_signal_19019) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_19022), .Q (new_AGEMA_signal_19023) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C (clk), .D (new_AGEMA_signal_19026), .Q (new_AGEMA_signal_19027) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_19030), .Q (new_AGEMA_signal_19031) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_19034), .Q (new_AGEMA_signal_19035) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C (clk), .D (new_AGEMA_signal_19038), .Q (new_AGEMA_signal_19039) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_19042), .Q (new_AGEMA_signal_19043) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C (clk), .D (new_AGEMA_signal_19046), .Q (new_AGEMA_signal_19047) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C (clk), .D (new_AGEMA_signal_19050), .Q (new_AGEMA_signal_19051) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_19054), .Q (new_AGEMA_signal_19055) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_19058), .Q (new_AGEMA_signal_19059) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C (clk), .D (new_AGEMA_signal_19062), .Q (new_AGEMA_signal_19063) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_19066), .Q (new_AGEMA_signal_19067) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_19070), .Q (new_AGEMA_signal_19071) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C (clk), .D (new_AGEMA_signal_19074), .Q (new_AGEMA_signal_19075) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_19078), .Q (new_AGEMA_signal_19079) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C (clk), .D (new_AGEMA_signal_19082), .Q (new_AGEMA_signal_19083) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C (clk), .D (new_AGEMA_signal_19086), .Q (new_AGEMA_signal_19087) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_19090), .Q (new_AGEMA_signal_19091) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_19094), .Q (new_AGEMA_signal_19095) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C (clk), .D (new_AGEMA_signal_19098), .Q (new_AGEMA_signal_19099) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_19102), .Q (new_AGEMA_signal_19103) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_19106), .Q (new_AGEMA_signal_19107) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C (clk), .D (new_AGEMA_signal_19110), .Q (new_AGEMA_signal_19111) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_19114), .Q (new_AGEMA_signal_19115) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C (clk), .D (new_AGEMA_signal_19118), .Q (new_AGEMA_signal_19119) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C (clk), .D (new_AGEMA_signal_19122), .Q (new_AGEMA_signal_19123) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_19126), .Q (new_AGEMA_signal_19127) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_19130), .Q (new_AGEMA_signal_19131) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C (clk), .D (new_AGEMA_signal_19134), .Q (new_AGEMA_signal_19135) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_19138), .Q (new_AGEMA_signal_19139) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_19142), .Q (new_AGEMA_signal_19143) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C (clk), .D (new_AGEMA_signal_19146), .Q (new_AGEMA_signal_19147) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_19150), .Q (new_AGEMA_signal_19151) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C (clk), .D (new_AGEMA_signal_19154), .Q (new_AGEMA_signal_19155) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C (clk), .D (new_AGEMA_signal_19158), .Q (new_AGEMA_signal_19159) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_19162), .Q (new_AGEMA_signal_19163) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_19166), .Q (new_AGEMA_signal_19167) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C (clk), .D (new_AGEMA_signal_19170), .Q (new_AGEMA_signal_19171) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_19174), .Q (new_AGEMA_signal_19175) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_19178), .Q (new_AGEMA_signal_19179) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C (clk), .D (new_AGEMA_signal_19182), .Q (new_AGEMA_signal_19183) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C (clk), .D (new_AGEMA_signal_19186), .Q (new_AGEMA_signal_19187) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_19190), .Q (new_AGEMA_signal_19191) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C (clk), .D (new_AGEMA_signal_19194), .Q (new_AGEMA_signal_19195) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_19198), .Q (new_AGEMA_signal_19199) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C (clk), .D (new_AGEMA_signal_19202), .Q (new_AGEMA_signal_19203) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C (clk), .D (new_AGEMA_signal_19206), .Q (new_AGEMA_signal_19207) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C (clk), .D (new_AGEMA_signal_19210), .Q (new_AGEMA_signal_19211) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_19214), .Q (new_AGEMA_signal_19215) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C (clk), .D (new_AGEMA_signal_19218), .Q (new_AGEMA_signal_19219) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_19222), .Q (new_AGEMA_signal_19223) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_19225), .Q (new_AGEMA_signal_19226) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C (clk), .D (new_AGEMA_signal_19228), .Q (new_AGEMA_signal_19229) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_19231), .Q (new_AGEMA_signal_19232) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_19234), .Q (new_AGEMA_signal_19235) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_19237), .Q (new_AGEMA_signal_19238) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C (clk), .D (new_AGEMA_signal_19240), .Q (new_AGEMA_signal_19241) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_19243), .Q (new_AGEMA_signal_19244) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_19246), .Q (new_AGEMA_signal_19247) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_19249), .Q (new_AGEMA_signal_19250) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C (clk), .D (new_AGEMA_signal_19252), .Q (new_AGEMA_signal_19253) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_19255), .Q (new_AGEMA_signal_19256) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_19258), .Q (new_AGEMA_signal_19259) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_19261), .Q (new_AGEMA_signal_19262) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C (clk), .D (new_AGEMA_signal_19264), .Q (new_AGEMA_signal_19265) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_19267), .Q (new_AGEMA_signal_19268) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_19270), .Q (new_AGEMA_signal_19271) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_19273), .Q (new_AGEMA_signal_19274) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C (clk), .D (new_AGEMA_signal_19276), .Q (new_AGEMA_signal_19277) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_19279), .Q (new_AGEMA_signal_19280) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_19282), .Q (new_AGEMA_signal_19283) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_19285), .Q (new_AGEMA_signal_19286) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C (clk), .D (new_AGEMA_signal_19288), .Q (new_AGEMA_signal_19289) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_19291), .Q (new_AGEMA_signal_19292) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_19294), .Q (new_AGEMA_signal_19295) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_19297), .Q (new_AGEMA_signal_19298) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C (clk), .D (new_AGEMA_signal_19300), .Q (new_AGEMA_signal_19301) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_19303), .Q (new_AGEMA_signal_19304) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_19306), .Q (new_AGEMA_signal_19307) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_19309), .Q (new_AGEMA_signal_19310) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C (clk), .D (new_AGEMA_signal_19312), .Q (new_AGEMA_signal_19313) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_19315), .Q (new_AGEMA_signal_19316) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_19318), .Q (new_AGEMA_signal_19319) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_19321), .Q (new_AGEMA_signal_19322) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C (clk), .D (new_AGEMA_signal_19324), .Q (new_AGEMA_signal_19325) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_19327), .Q (new_AGEMA_signal_19328) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_19330), .Q (new_AGEMA_signal_19331) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_19333), .Q (new_AGEMA_signal_19334) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C (clk), .D (new_AGEMA_signal_19336), .Q (new_AGEMA_signal_19337) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_19339), .Q (new_AGEMA_signal_19340) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_19342), .Q (new_AGEMA_signal_19343) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_19345), .Q (new_AGEMA_signal_19346) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C (clk), .D (new_AGEMA_signal_19348), .Q (new_AGEMA_signal_19349) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_19351), .Q (new_AGEMA_signal_19352) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_19354), .Q (new_AGEMA_signal_19355) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_19357), .Q (new_AGEMA_signal_19358) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C (clk), .D (new_AGEMA_signal_19360), .Q (new_AGEMA_signal_19361) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_19363), .Q (new_AGEMA_signal_19364) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_19366), .Q (new_AGEMA_signal_19367) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_19369), .Q (new_AGEMA_signal_19370) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C (clk), .D (new_AGEMA_signal_19372), .Q (new_AGEMA_signal_19373) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_19375), .Q (new_AGEMA_signal_19376) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_19378), .Q (new_AGEMA_signal_19379) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_19381), .Q (new_AGEMA_signal_19382) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C (clk), .D (new_AGEMA_signal_19384), .Q (new_AGEMA_signal_19385) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_19387), .Q (new_AGEMA_signal_19388) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_19390), .Q (new_AGEMA_signal_19391) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_19393), .Q (new_AGEMA_signal_19394) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C (clk), .D (new_AGEMA_signal_19396), .Q (new_AGEMA_signal_19397) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_19399), .Q (new_AGEMA_signal_19400) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_19402), .Q (new_AGEMA_signal_19403) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_19405), .Q (new_AGEMA_signal_19406) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C (clk), .D (new_AGEMA_signal_19408), .Q (new_AGEMA_signal_19409) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C (clk), .D (new_AGEMA_signal_19411), .Q (new_AGEMA_signal_19412) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C (clk), .D (new_AGEMA_signal_19414), .Q (new_AGEMA_signal_19415) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C (clk), .D (new_AGEMA_signal_19417), .Q (new_AGEMA_signal_19418) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C (clk), .D (new_AGEMA_signal_19420), .Q (new_AGEMA_signal_19421) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C (clk), .D (new_AGEMA_signal_19423), .Q (new_AGEMA_signal_19424) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C (clk), .D (new_AGEMA_signal_19426), .Q (new_AGEMA_signal_19427) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C (clk), .D (new_AGEMA_signal_19429), .Q (new_AGEMA_signal_19430) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C (clk), .D (new_AGEMA_signal_19432), .Q (new_AGEMA_signal_19433) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C (clk), .D (new_AGEMA_signal_19435), .Q (new_AGEMA_signal_19436) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C (clk), .D (new_AGEMA_signal_19438), .Q (new_AGEMA_signal_19439) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C (clk), .D (new_AGEMA_signal_19441), .Q (new_AGEMA_signal_19442) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C (clk), .D (new_AGEMA_signal_19444), .Q (new_AGEMA_signal_19445) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C (clk), .D (new_AGEMA_signal_19447), .Q (new_AGEMA_signal_19448) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C (clk), .D (new_AGEMA_signal_19450), .Q (new_AGEMA_signal_19451) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C (clk), .D (new_AGEMA_signal_19453), .Q (new_AGEMA_signal_19454) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C (clk), .D (new_AGEMA_signal_19456), .Q (new_AGEMA_signal_19457) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C (clk), .D (new_AGEMA_signal_19459), .Q (new_AGEMA_signal_19460) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C (clk), .D (new_AGEMA_signal_19462), .Q (new_AGEMA_signal_19463) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C (clk), .D (new_AGEMA_signal_19465), .Q (new_AGEMA_signal_19466) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C (clk), .D (new_AGEMA_signal_19468), .Q (new_AGEMA_signal_19469) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C (clk), .D (new_AGEMA_signal_19471), .Q (new_AGEMA_signal_19472) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C (clk), .D (new_AGEMA_signal_19474), .Q (new_AGEMA_signal_19475) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C (clk), .D (new_AGEMA_signal_19477), .Q (new_AGEMA_signal_19478) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C (clk), .D (new_AGEMA_signal_19480), .Q (new_AGEMA_signal_19481) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C (clk), .D (new_AGEMA_signal_19483), .Q (new_AGEMA_signal_19484) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C (clk), .D (new_AGEMA_signal_19486), .Q (new_AGEMA_signal_19487) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C (clk), .D (new_AGEMA_signal_19489), .Q (new_AGEMA_signal_19490) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C (clk), .D (new_AGEMA_signal_19492), .Q (new_AGEMA_signal_19493) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C (clk), .D (new_AGEMA_signal_19495), .Q (new_AGEMA_signal_19496) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C (clk), .D (new_AGEMA_signal_19498), .Q (new_AGEMA_signal_19499) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C (clk), .D (new_AGEMA_signal_19501), .Q (new_AGEMA_signal_19502) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C (clk), .D (new_AGEMA_signal_19504), .Q (new_AGEMA_signal_19505) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C (clk), .D (new_AGEMA_signal_19507), .Q (new_AGEMA_signal_19508) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C (clk), .D (new_AGEMA_signal_19510), .Q (new_AGEMA_signal_19511) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C (clk), .D (new_AGEMA_signal_19513), .Q (new_AGEMA_signal_19514) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C (clk), .D (new_AGEMA_signal_19516), .Q (new_AGEMA_signal_19517) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C (clk), .D (new_AGEMA_signal_19519), .Q (new_AGEMA_signal_19520) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C (clk), .D (new_AGEMA_signal_19522), .Q (new_AGEMA_signal_19523) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C (clk), .D (new_AGEMA_signal_19525), .Q (new_AGEMA_signal_19526) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C (clk), .D (new_AGEMA_signal_19528), .Q (new_AGEMA_signal_19529) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C (clk), .D (new_AGEMA_signal_19531), .Q (new_AGEMA_signal_19532) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C (clk), .D (new_AGEMA_signal_19534), .Q (new_AGEMA_signal_19535) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C (clk), .D (new_AGEMA_signal_19537), .Q (new_AGEMA_signal_19538) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C (clk), .D (new_AGEMA_signal_19540), .Q (new_AGEMA_signal_19541) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C (clk), .D (new_AGEMA_signal_19543), .Q (new_AGEMA_signal_19544) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C (clk), .D (new_AGEMA_signal_19546), .Q (new_AGEMA_signal_19547) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C (clk), .D (new_AGEMA_signal_19549), .Q (new_AGEMA_signal_19550) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C (clk), .D (new_AGEMA_signal_19552), .Q (new_AGEMA_signal_19553) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C (clk), .D (new_AGEMA_signal_19555), .Q (new_AGEMA_signal_19556) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C (clk), .D (new_AGEMA_signal_19558), .Q (new_AGEMA_signal_19559) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C (clk), .D (new_AGEMA_signal_19561), .Q (new_AGEMA_signal_19562) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C (clk), .D (new_AGEMA_signal_19564), .Q (new_AGEMA_signal_19565) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C (clk), .D (new_AGEMA_signal_19567), .Q (new_AGEMA_signal_19568) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C (clk), .D (new_AGEMA_signal_19570), .Q (new_AGEMA_signal_19571) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C (clk), .D (new_AGEMA_signal_19573), .Q (new_AGEMA_signal_19574) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C (clk), .D (new_AGEMA_signal_19576), .Q (new_AGEMA_signal_19577) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C (clk), .D (new_AGEMA_signal_19579), .Q (new_AGEMA_signal_19580) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C (clk), .D (new_AGEMA_signal_19582), .Q (new_AGEMA_signal_19583) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C (clk), .D (new_AGEMA_signal_19585), .Q (new_AGEMA_signal_19586) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C (clk), .D (new_AGEMA_signal_19588), .Q (new_AGEMA_signal_19589) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C (clk), .D (new_AGEMA_signal_19591), .Q (new_AGEMA_signal_19592) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C (clk), .D (new_AGEMA_signal_19594), .Q (new_AGEMA_signal_19595) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C (clk), .D (new_AGEMA_signal_19597), .Q (new_AGEMA_signal_19598) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C (clk), .D (new_AGEMA_signal_19600), .Q (new_AGEMA_signal_19601) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C (clk), .D (new_AGEMA_signal_19603), .Q (new_AGEMA_signal_19604) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C (clk), .D (new_AGEMA_signal_19606), .Q (new_AGEMA_signal_19607) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C (clk), .D (new_AGEMA_signal_19609), .Q (new_AGEMA_signal_19610) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C (clk), .D (new_AGEMA_signal_19612), .Q (new_AGEMA_signal_19613) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C (clk), .D (new_AGEMA_signal_19615), .Q (new_AGEMA_signal_19616) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C (clk), .D (new_AGEMA_signal_19618), .Q (new_AGEMA_signal_19619) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C (clk), .D (new_AGEMA_signal_19621), .Q (new_AGEMA_signal_19622) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C (clk), .D (new_AGEMA_signal_19624), .Q (new_AGEMA_signal_19625) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C (clk), .D (new_AGEMA_signal_19627), .Q (new_AGEMA_signal_19628) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C (clk), .D (new_AGEMA_signal_19630), .Q (new_AGEMA_signal_19631) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C (clk), .D (new_AGEMA_signal_19633), .Q (new_AGEMA_signal_19634) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C (clk), .D (new_AGEMA_signal_19636), .Q (new_AGEMA_signal_19637) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C (clk), .D (new_AGEMA_signal_19639), .Q (new_AGEMA_signal_19640) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C (clk), .D (new_AGEMA_signal_19642), .Q (new_AGEMA_signal_19643) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C (clk), .D (new_AGEMA_signal_19645), .Q (new_AGEMA_signal_19646) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C (clk), .D (new_AGEMA_signal_19648), .Q (new_AGEMA_signal_19649) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C (clk), .D (new_AGEMA_signal_19651), .Q (new_AGEMA_signal_19652) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C (clk), .D (new_AGEMA_signal_19654), .Q (new_AGEMA_signal_19655) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C (clk), .D (new_AGEMA_signal_19657), .Q (new_AGEMA_signal_19658) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C (clk), .D (new_AGEMA_signal_19660), .Q (new_AGEMA_signal_19661) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C (clk), .D (new_AGEMA_signal_19663), .Q (new_AGEMA_signal_19664) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C (clk), .D (new_AGEMA_signal_19666), .Q (new_AGEMA_signal_19667) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C (clk), .D (new_AGEMA_signal_19669), .Q (new_AGEMA_signal_19670) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C (clk), .D (new_AGEMA_signal_19672), .Q (new_AGEMA_signal_19673) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C (clk), .D (new_AGEMA_signal_19675), .Q (new_AGEMA_signal_19676) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C (clk), .D (new_AGEMA_signal_19678), .Q (new_AGEMA_signal_19679) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C (clk), .D (new_AGEMA_signal_19681), .Q (new_AGEMA_signal_19682) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C (clk), .D (new_AGEMA_signal_19684), .Q (new_AGEMA_signal_19685) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C (clk), .D (new_AGEMA_signal_19687), .Q (new_AGEMA_signal_19688) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C (clk), .D (new_AGEMA_signal_19690), .Q (new_AGEMA_signal_19691) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C (clk), .D (new_AGEMA_signal_19693), .Q (new_AGEMA_signal_19694) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C (clk), .D (new_AGEMA_signal_19696), .Q (new_AGEMA_signal_19697) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C (clk), .D (new_AGEMA_signal_19699), .Q (new_AGEMA_signal_19700) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C (clk), .D (new_AGEMA_signal_19702), .Q (new_AGEMA_signal_19703) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C (clk), .D (new_AGEMA_signal_19705), .Q (new_AGEMA_signal_19706) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C (clk), .D (new_AGEMA_signal_19708), .Q (new_AGEMA_signal_19709) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C (clk), .D (new_AGEMA_signal_19711), .Q (new_AGEMA_signal_19712) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C (clk), .D (new_AGEMA_signal_19714), .Q (new_AGEMA_signal_19715) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C (clk), .D (new_AGEMA_signal_19717), .Q (new_AGEMA_signal_19718) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C (clk), .D (new_AGEMA_signal_19720), .Q (new_AGEMA_signal_19721) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C (clk), .D (new_AGEMA_signal_19723), .Q (new_AGEMA_signal_19724) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C (clk), .D (new_AGEMA_signal_19726), .Q (new_AGEMA_signal_19727) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C (clk), .D (new_AGEMA_signal_19729), .Q (new_AGEMA_signal_19730) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C (clk), .D (new_AGEMA_signal_19732), .Q (new_AGEMA_signal_19733) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C (clk), .D (new_AGEMA_signal_19735), .Q (new_AGEMA_signal_19736) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C (clk), .D (new_AGEMA_signal_19738), .Q (new_AGEMA_signal_19739) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C (clk), .D (new_AGEMA_signal_19741), .Q (new_AGEMA_signal_19742) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C (clk), .D (new_AGEMA_signal_19744), .Q (new_AGEMA_signal_19745) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C (clk), .D (new_AGEMA_signal_19747), .Q (new_AGEMA_signal_19748) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C (clk), .D (new_AGEMA_signal_19750), .Q (new_AGEMA_signal_19751) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C (clk), .D (new_AGEMA_signal_19753), .Q (new_AGEMA_signal_19754) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C (clk), .D (new_AGEMA_signal_19756), .Q (new_AGEMA_signal_19757) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C (clk), .D (new_AGEMA_signal_19759), .Q (new_AGEMA_signal_19760) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C (clk), .D (new_AGEMA_signal_19762), .Q (new_AGEMA_signal_19763) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C (clk), .D (new_AGEMA_signal_19765), .Q (new_AGEMA_signal_19766) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C (clk), .D (new_AGEMA_signal_19768), .Q (new_AGEMA_signal_19769) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C (clk), .D (new_AGEMA_signal_19771), .Q (new_AGEMA_signal_19772) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C (clk), .D (new_AGEMA_signal_19774), .Q (new_AGEMA_signal_19775) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C (clk), .D (new_AGEMA_signal_19777), .Q (new_AGEMA_signal_19778) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C (clk), .D (new_AGEMA_signal_19780), .Q (new_AGEMA_signal_19781) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C (clk), .D (new_AGEMA_signal_19783), .Q (new_AGEMA_signal_19784) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C (clk), .D (new_AGEMA_signal_19786), .Q (new_AGEMA_signal_19787) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C (clk), .D (new_AGEMA_signal_19789), .Q (new_AGEMA_signal_19790) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C (clk), .D (new_AGEMA_signal_19792), .Q (new_AGEMA_signal_19793) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C (clk), .D (new_AGEMA_signal_19795), .Q (new_AGEMA_signal_19796) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C (clk), .D (new_AGEMA_signal_19798), .Q (new_AGEMA_signal_19799) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C (clk), .D (new_AGEMA_signal_19801), .Q (new_AGEMA_signal_19802) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C (clk), .D (new_AGEMA_signal_19804), .Q (new_AGEMA_signal_19805) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C (clk), .D (new_AGEMA_signal_19807), .Q (new_AGEMA_signal_19808) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C (clk), .D (new_AGEMA_signal_19810), .Q (new_AGEMA_signal_19811) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C (clk), .D (new_AGEMA_signal_19813), .Q (new_AGEMA_signal_19814) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C (clk), .D (new_AGEMA_signal_19816), .Q (new_AGEMA_signal_19817) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C (clk), .D (new_AGEMA_signal_19819), .Q (new_AGEMA_signal_19820) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C (clk), .D (new_AGEMA_signal_19822), .Q (new_AGEMA_signal_19823) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C (clk), .D (new_AGEMA_signal_19825), .Q (new_AGEMA_signal_19826) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C (clk), .D (new_AGEMA_signal_19828), .Q (new_AGEMA_signal_19829) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C (clk), .D (new_AGEMA_signal_19831), .Q (new_AGEMA_signal_19832) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C (clk), .D (new_AGEMA_signal_19834), .Q (new_AGEMA_signal_19835) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C (clk), .D (new_AGEMA_signal_19837), .Q (new_AGEMA_signal_19838) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C (clk), .D (new_AGEMA_signal_19840), .Q (new_AGEMA_signal_19841) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C (clk), .D (new_AGEMA_signal_19843), .Q (new_AGEMA_signal_19844) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C (clk), .D (new_AGEMA_signal_19846), .Q (new_AGEMA_signal_19847) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C (clk), .D (new_AGEMA_signal_19849), .Q (new_AGEMA_signal_19850) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C (clk), .D (new_AGEMA_signal_19852), .Q (new_AGEMA_signal_19853) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C (clk), .D (new_AGEMA_signal_19855), .Q (new_AGEMA_signal_19856) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C (clk), .D (new_AGEMA_signal_19858), .Q (new_AGEMA_signal_19859) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C (clk), .D (new_AGEMA_signal_19861), .Q (new_AGEMA_signal_19862) ) ;
    buf_clk new_AGEMA_reg_buffer_7141 ( .C (clk), .D (new_AGEMA_signal_19864), .Q (new_AGEMA_signal_19865) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C (clk), .D (new_AGEMA_signal_19867), .Q (new_AGEMA_signal_19868) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C (clk), .D (new_AGEMA_signal_19870), .Q (new_AGEMA_signal_19871) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C (clk), .D (new_AGEMA_signal_19873), .Q (new_AGEMA_signal_19874) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C (clk), .D (new_AGEMA_signal_19876), .Q (new_AGEMA_signal_19877) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C (clk), .D (new_AGEMA_signal_19879), .Q (new_AGEMA_signal_19880) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C (clk), .D (new_AGEMA_signal_19882), .Q (new_AGEMA_signal_19883) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C (clk), .D (new_AGEMA_signal_19885), .Q (new_AGEMA_signal_19886) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C (clk), .D (new_AGEMA_signal_19888), .Q (new_AGEMA_signal_19889) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C (clk), .D (new_AGEMA_signal_19891), .Q (new_AGEMA_signal_19892) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C (clk), .D (new_AGEMA_signal_19894), .Q (new_AGEMA_signal_19895) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C (clk), .D (new_AGEMA_signal_19897), .Q (new_AGEMA_signal_19898) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C (clk), .D (new_AGEMA_signal_19900), .Q (new_AGEMA_signal_19901) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C (clk), .D (new_AGEMA_signal_19903), .Q (new_AGEMA_signal_19904) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C (clk), .D (new_AGEMA_signal_19906), .Q (new_AGEMA_signal_19907) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C (clk), .D (new_AGEMA_signal_19909), .Q (new_AGEMA_signal_19910) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C (clk), .D (new_AGEMA_signal_19912), .Q (new_AGEMA_signal_19913) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C (clk), .D (new_AGEMA_signal_19915), .Q (new_AGEMA_signal_19916) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C (clk), .D (new_AGEMA_signal_19918), .Q (new_AGEMA_signal_19919) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C (clk), .D (new_AGEMA_signal_19921), .Q (new_AGEMA_signal_19922) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C (clk), .D (new_AGEMA_signal_19924), .Q (new_AGEMA_signal_19925) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C (clk), .D (new_AGEMA_signal_19927), .Q (new_AGEMA_signal_19928) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C (clk), .D (new_AGEMA_signal_19930), .Q (new_AGEMA_signal_19931) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C (clk), .D (new_AGEMA_signal_19933), .Q (new_AGEMA_signal_19934) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C (clk), .D (new_AGEMA_signal_19936), .Q (new_AGEMA_signal_19937) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C (clk), .D (new_AGEMA_signal_19939), .Q (new_AGEMA_signal_19940) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C (clk), .D (new_AGEMA_signal_19942), .Q (new_AGEMA_signal_19943) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C (clk), .D (new_AGEMA_signal_19945), .Q (new_AGEMA_signal_19946) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C (clk), .D (new_AGEMA_signal_19948), .Q (new_AGEMA_signal_19949) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C (clk), .D (new_AGEMA_signal_19951), .Q (new_AGEMA_signal_19952) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C (clk), .D (new_AGEMA_signal_19954), .Q (new_AGEMA_signal_19955) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C (clk), .D (new_AGEMA_signal_19957), .Q (new_AGEMA_signal_19958) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C (clk), .D (new_AGEMA_signal_19960), .Q (new_AGEMA_signal_19961) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C (clk), .D (new_AGEMA_signal_19963), .Q (new_AGEMA_signal_19964) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C (clk), .D (new_AGEMA_signal_19966), .Q (new_AGEMA_signal_19967) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C (clk), .D (new_AGEMA_signal_19969), .Q (new_AGEMA_signal_19970) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C (clk), .D (new_AGEMA_signal_19972), .Q (new_AGEMA_signal_19973) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C (clk), .D (new_AGEMA_signal_19975), .Q (new_AGEMA_signal_19976) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C (clk), .D (new_AGEMA_signal_19978), .Q (new_AGEMA_signal_19979) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C (clk), .D (new_AGEMA_signal_19981), .Q (new_AGEMA_signal_19982) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C (clk), .D (new_AGEMA_signal_19984), .Q (new_AGEMA_signal_19985) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C (clk), .D (new_AGEMA_signal_19987), .Q (new_AGEMA_signal_19988) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C (clk), .D (new_AGEMA_signal_19990), .Q (new_AGEMA_signal_19991) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C (clk), .D (new_AGEMA_signal_19993), .Q (new_AGEMA_signal_19994) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C (clk), .D (new_AGEMA_signal_19996), .Q (new_AGEMA_signal_19997) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C (clk), .D (new_AGEMA_signal_19999), .Q (new_AGEMA_signal_20000) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C (clk), .D (new_AGEMA_signal_20002), .Q (new_AGEMA_signal_20003) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C (clk), .D (new_AGEMA_signal_20005), .Q (new_AGEMA_signal_20006) ) ;
    buf_clk new_AGEMA_reg_buffer_7285 ( .C (clk), .D (new_AGEMA_signal_20008), .Q (new_AGEMA_signal_20009) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C (clk), .D (new_AGEMA_signal_20011), .Q (new_AGEMA_signal_20012) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C (clk), .D (new_AGEMA_signal_20014), .Q (new_AGEMA_signal_20015) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C (clk), .D (new_AGEMA_signal_20017), .Q (new_AGEMA_signal_20018) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C (clk), .D (new_AGEMA_signal_20020), .Q (new_AGEMA_signal_20021) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C (clk), .D (new_AGEMA_signal_20023), .Q (new_AGEMA_signal_20024) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C (clk), .D (new_AGEMA_signal_20026), .Q (new_AGEMA_signal_20027) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C (clk), .D (new_AGEMA_signal_20029), .Q (new_AGEMA_signal_20030) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C (clk), .D (new_AGEMA_signal_20032), .Q (new_AGEMA_signal_20033) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C (clk), .D (new_AGEMA_signal_20035), .Q (new_AGEMA_signal_20036) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C (clk), .D (new_AGEMA_signal_20038), .Q (new_AGEMA_signal_20039) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C (clk), .D (new_AGEMA_signal_20041), .Q (new_AGEMA_signal_20042) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C (clk), .D (new_AGEMA_signal_20044), .Q (new_AGEMA_signal_20045) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C (clk), .D (new_AGEMA_signal_20047), .Q (new_AGEMA_signal_20048) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C (clk), .D (new_AGEMA_signal_20050), .Q (new_AGEMA_signal_20051) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C (clk), .D (new_AGEMA_signal_20053), .Q (new_AGEMA_signal_20054) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C (clk), .D (new_AGEMA_signal_20056), .Q (new_AGEMA_signal_20057) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C (clk), .D (new_AGEMA_signal_20059), .Q (new_AGEMA_signal_20060) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C (clk), .D (new_AGEMA_signal_20062), .Q (new_AGEMA_signal_20063) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C (clk), .D (new_AGEMA_signal_20065), .Q (new_AGEMA_signal_20066) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C (clk), .D (new_AGEMA_signal_20068), .Q (new_AGEMA_signal_20069) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C (clk), .D (new_AGEMA_signal_20071), .Q (new_AGEMA_signal_20072) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C (clk), .D (new_AGEMA_signal_20074), .Q (new_AGEMA_signal_20075) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C (clk), .D (new_AGEMA_signal_20077), .Q (new_AGEMA_signal_20078) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C (clk), .D (new_AGEMA_signal_20080), .Q (new_AGEMA_signal_20081) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C (clk), .D (new_AGEMA_signal_20083), .Q (new_AGEMA_signal_20084) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C (clk), .D (new_AGEMA_signal_20086), .Q (new_AGEMA_signal_20087) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C (clk), .D (new_AGEMA_signal_20089), .Q (new_AGEMA_signal_20090) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C (clk), .D (new_AGEMA_signal_20092), .Q (new_AGEMA_signal_20093) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C (clk), .D (new_AGEMA_signal_20095), .Q (new_AGEMA_signal_20096) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C (clk), .D (new_AGEMA_signal_20098), .Q (new_AGEMA_signal_20099) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C (clk), .D (new_AGEMA_signal_20101), .Q (new_AGEMA_signal_20102) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C (clk), .D (new_AGEMA_signal_20104), .Q (new_AGEMA_signal_20105) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C (clk), .D (new_AGEMA_signal_20107), .Q (new_AGEMA_signal_20108) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C (clk), .D (new_AGEMA_signal_20110), .Q (new_AGEMA_signal_20111) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C (clk), .D (new_AGEMA_signal_20113), .Q (new_AGEMA_signal_20114) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C (clk), .D (new_AGEMA_signal_20116), .Q (new_AGEMA_signal_20117) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C (clk), .D (new_AGEMA_signal_20119), .Q (new_AGEMA_signal_20120) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C (clk), .D (new_AGEMA_signal_20122), .Q (new_AGEMA_signal_20123) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C (clk), .D (new_AGEMA_signal_20125), .Q (new_AGEMA_signal_20126) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C (clk), .D (new_AGEMA_signal_20128), .Q (new_AGEMA_signal_20129) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C (clk), .D (new_AGEMA_signal_20131), .Q (new_AGEMA_signal_20132) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C (clk), .D (new_AGEMA_signal_20134), .Q (new_AGEMA_signal_20135) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C (clk), .D (new_AGEMA_signal_20137), .Q (new_AGEMA_signal_20138) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C (clk), .D (new_AGEMA_signal_20140), .Q (new_AGEMA_signal_20141) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C (clk), .D (new_AGEMA_signal_20143), .Q (new_AGEMA_signal_20144) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C (clk), .D (new_AGEMA_signal_20146), .Q (new_AGEMA_signal_20147) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C (clk), .D (new_AGEMA_signal_20149), .Q (new_AGEMA_signal_20150) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C (clk), .D (new_AGEMA_signal_20152), .Q (new_AGEMA_signal_20153) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C (clk), .D (new_AGEMA_signal_20155), .Q (new_AGEMA_signal_20156) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C (clk), .D (new_AGEMA_signal_20158), .Q (new_AGEMA_signal_20159) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C (clk), .D (new_AGEMA_signal_20161), .Q (new_AGEMA_signal_20162) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C (clk), .D (new_AGEMA_signal_20164), .Q (new_AGEMA_signal_20165) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C (clk), .D (new_AGEMA_signal_20167), .Q (new_AGEMA_signal_20168) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C (clk), .D (new_AGEMA_signal_20170), .Q (new_AGEMA_signal_20171) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C (clk), .D (new_AGEMA_signal_20173), .Q (new_AGEMA_signal_20174) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C (clk), .D (new_AGEMA_signal_20176), .Q (new_AGEMA_signal_20177) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C (clk), .D (new_AGEMA_signal_20179), .Q (new_AGEMA_signal_20180) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C (clk), .D (new_AGEMA_signal_20182), .Q (new_AGEMA_signal_20183) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C (clk), .D (new_AGEMA_signal_20185), .Q (new_AGEMA_signal_20186) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C (clk), .D (new_AGEMA_signal_20188), .Q (new_AGEMA_signal_20189) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C (clk), .D (new_AGEMA_signal_20191), .Q (new_AGEMA_signal_20192) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C (clk), .D (new_AGEMA_signal_20194), .Q (new_AGEMA_signal_20195) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C (clk), .D (new_AGEMA_signal_20197), .Q (new_AGEMA_signal_20198) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C (clk), .D (new_AGEMA_signal_20200), .Q (new_AGEMA_signal_20201) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C (clk), .D (new_AGEMA_signal_20203), .Q (new_AGEMA_signal_20204) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C (clk), .D (new_AGEMA_signal_20206), .Q (new_AGEMA_signal_20207) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C (clk), .D (new_AGEMA_signal_20209), .Q (new_AGEMA_signal_20210) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C (clk), .D (new_AGEMA_signal_20212), .Q (new_AGEMA_signal_20213) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C (clk), .D (new_AGEMA_signal_20215), .Q (new_AGEMA_signal_20216) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C (clk), .D (new_AGEMA_signal_20218), .Q (new_AGEMA_signal_20219) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C (clk), .D (new_AGEMA_signal_20221), .Q (new_AGEMA_signal_20222) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C (clk), .D (new_AGEMA_signal_20224), .Q (new_AGEMA_signal_20225) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C (clk), .D (new_AGEMA_signal_20227), .Q (new_AGEMA_signal_20228) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C (clk), .D (new_AGEMA_signal_20230), .Q (new_AGEMA_signal_20231) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C (clk), .D (new_AGEMA_signal_20233), .Q (new_AGEMA_signal_20234) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C (clk), .D (new_AGEMA_signal_20236), .Q (new_AGEMA_signal_20237) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C (clk), .D (new_AGEMA_signal_20239), .Q (new_AGEMA_signal_20240) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C (clk), .D (new_AGEMA_signal_20242), .Q (new_AGEMA_signal_20243) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C (clk), .D (new_AGEMA_signal_20245), .Q (new_AGEMA_signal_20246) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C (clk), .D (new_AGEMA_signal_20248), .Q (new_AGEMA_signal_20249) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C (clk), .D (new_AGEMA_signal_20251), .Q (new_AGEMA_signal_20252) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C (clk), .D (new_AGEMA_signal_20254), .Q (new_AGEMA_signal_20255) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C (clk), .D (new_AGEMA_signal_20257), .Q (new_AGEMA_signal_20258) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C (clk), .D (new_AGEMA_signal_20260), .Q (new_AGEMA_signal_20261) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C (clk), .D (new_AGEMA_signal_20263), .Q (new_AGEMA_signal_20264) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C (clk), .D (new_AGEMA_signal_20266), .Q (new_AGEMA_signal_20267) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C (clk), .D (new_AGEMA_signal_20269), .Q (new_AGEMA_signal_20270) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C (clk), .D (new_AGEMA_signal_20272), .Q (new_AGEMA_signal_20273) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C (clk), .D (new_AGEMA_signal_20275), .Q (new_AGEMA_signal_20276) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C (clk), .D (new_AGEMA_signal_20278), .Q (new_AGEMA_signal_20279) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C (clk), .D (new_AGEMA_signal_20281), .Q (new_AGEMA_signal_20282) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C (clk), .D (new_AGEMA_signal_20284), .Q (new_AGEMA_signal_20285) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C (clk), .D (new_AGEMA_signal_20287), .Q (new_AGEMA_signal_20288) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C (clk), .D (new_AGEMA_signal_20290), .Q (new_AGEMA_signal_20291) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C (clk), .D (new_AGEMA_signal_20293), .Q (new_AGEMA_signal_20294) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C (clk), .D (new_AGEMA_signal_20296), .Q (new_AGEMA_signal_20297) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C (clk), .D (new_AGEMA_signal_20299), .Q (new_AGEMA_signal_20300) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C (clk), .D (new_AGEMA_signal_20302), .Q (new_AGEMA_signal_20303) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C (clk), .D (new_AGEMA_signal_20305), .Q (new_AGEMA_signal_20306) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C (clk), .D (new_AGEMA_signal_20308), .Q (new_AGEMA_signal_20309) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C (clk), .D (new_AGEMA_signal_20311), .Q (new_AGEMA_signal_20312) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C (clk), .D (new_AGEMA_signal_20314), .Q (new_AGEMA_signal_20315) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C (clk), .D (new_AGEMA_signal_20317), .Q (new_AGEMA_signal_20318) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C (clk), .D (new_AGEMA_signal_20320), .Q (new_AGEMA_signal_20321) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C (clk), .D (new_AGEMA_signal_20323), .Q (new_AGEMA_signal_20324) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C (clk), .D (new_AGEMA_signal_20326), .Q (new_AGEMA_signal_20327) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C (clk), .D (new_AGEMA_signal_20329), .Q (new_AGEMA_signal_20330) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C (clk), .D (new_AGEMA_signal_20332), .Q (new_AGEMA_signal_20333) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C (clk), .D (new_AGEMA_signal_20335), .Q (new_AGEMA_signal_20336) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C (clk), .D (new_AGEMA_signal_20338), .Q (new_AGEMA_signal_20339) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C (clk), .D (new_AGEMA_signal_20341), .Q (new_AGEMA_signal_20342) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C (clk), .D (new_AGEMA_signal_20344), .Q (new_AGEMA_signal_20345) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C (clk), .D (new_AGEMA_signal_20347), .Q (new_AGEMA_signal_20348) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C (clk), .D (new_AGEMA_signal_20350), .Q (new_AGEMA_signal_20351) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C (clk), .D (new_AGEMA_signal_20353), .Q (new_AGEMA_signal_20354) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C (clk), .D (new_AGEMA_signal_20356), .Q (new_AGEMA_signal_20357) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C (clk), .D (new_AGEMA_signal_20359), .Q (new_AGEMA_signal_20360) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C (clk), .D (new_AGEMA_signal_20362), .Q (new_AGEMA_signal_20363) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C (clk), .D (new_AGEMA_signal_20365), .Q (new_AGEMA_signal_20366) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C (clk), .D (new_AGEMA_signal_20368), .Q (new_AGEMA_signal_20369) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C (clk), .D (new_AGEMA_signal_20371), .Q (new_AGEMA_signal_20372) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C (clk), .D (new_AGEMA_signal_20374), .Q (new_AGEMA_signal_20375) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C (clk), .D (new_AGEMA_signal_20377), .Q (new_AGEMA_signal_20378) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C (clk), .D (new_AGEMA_signal_20380), .Q (new_AGEMA_signal_20381) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C (clk), .D (new_AGEMA_signal_20383), .Q (new_AGEMA_signal_20384) ) ;
    buf_clk new_AGEMA_reg_buffer_7663 ( .C (clk), .D (new_AGEMA_signal_20386), .Q (new_AGEMA_signal_20387) ) ;
    buf_clk new_AGEMA_reg_buffer_7666 ( .C (clk), .D (new_AGEMA_signal_20389), .Q (new_AGEMA_signal_20390) ) ;
    buf_clk new_AGEMA_reg_buffer_7669 ( .C (clk), .D (new_AGEMA_signal_20392), .Q (new_AGEMA_signal_20393) ) ;
    buf_clk new_AGEMA_reg_buffer_7672 ( .C (clk), .D (new_AGEMA_signal_20395), .Q (new_AGEMA_signal_20396) ) ;
    buf_clk new_AGEMA_reg_buffer_7675 ( .C (clk), .D (new_AGEMA_signal_20398), .Q (new_AGEMA_signal_20399) ) ;
    buf_clk new_AGEMA_reg_buffer_7678 ( .C (clk), .D (new_AGEMA_signal_20401), .Q (new_AGEMA_signal_20402) ) ;
    buf_clk new_AGEMA_reg_buffer_7681 ( .C (clk), .D (new_AGEMA_signal_20404), .Q (new_AGEMA_signal_20405) ) ;
    buf_clk new_AGEMA_reg_buffer_7684 ( .C (clk), .D (new_AGEMA_signal_20407), .Q (new_AGEMA_signal_20408) ) ;
    buf_clk new_AGEMA_reg_buffer_7687 ( .C (clk), .D (new_AGEMA_signal_20410), .Q (new_AGEMA_signal_20411) ) ;
    buf_clk new_AGEMA_reg_buffer_7690 ( .C (clk), .D (new_AGEMA_signal_20413), .Q (new_AGEMA_signal_20414) ) ;
    buf_clk new_AGEMA_reg_buffer_7693 ( .C (clk), .D (new_AGEMA_signal_20416), .Q (new_AGEMA_signal_20417) ) ;
    buf_clk new_AGEMA_reg_buffer_7696 ( .C (clk), .D (new_AGEMA_signal_20419), .Q (new_AGEMA_signal_20420) ) ;
    buf_clk new_AGEMA_reg_buffer_7699 ( .C (clk), .D (new_AGEMA_signal_20422), .Q (new_AGEMA_signal_20423) ) ;
    buf_clk new_AGEMA_reg_buffer_7702 ( .C (clk), .D (new_AGEMA_signal_20425), .Q (new_AGEMA_signal_20426) ) ;
    buf_clk new_AGEMA_reg_buffer_7705 ( .C (clk), .D (new_AGEMA_signal_20428), .Q (new_AGEMA_signal_20429) ) ;
    buf_clk new_AGEMA_reg_buffer_7708 ( .C (clk), .D (new_AGEMA_signal_20431), .Q (new_AGEMA_signal_20432) ) ;
    buf_clk new_AGEMA_reg_buffer_7711 ( .C (clk), .D (new_AGEMA_signal_20434), .Q (new_AGEMA_signal_20435) ) ;
    buf_clk new_AGEMA_reg_buffer_7714 ( .C (clk), .D (new_AGEMA_signal_20437), .Q (new_AGEMA_signal_20438) ) ;
    buf_clk new_AGEMA_reg_buffer_7717 ( .C (clk), .D (new_AGEMA_signal_20440), .Q (new_AGEMA_signal_20441) ) ;
    buf_clk new_AGEMA_reg_buffer_7720 ( .C (clk), .D (new_AGEMA_signal_20443), .Q (new_AGEMA_signal_20444) ) ;
    buf_clk new_AGEMA_reg_buffer_7723 ( .C (clk), .D (new_AGEMA_signal_20446), .Q (new_AGEMA_signal_20447) ) ;
    buf_clk new_AGEMA_reg_buffer_7726 ( .C (clk), .D (new_AGEMA_signal_20449), .Q (new_AGEMA_signal_20450) ) ;
    buf_clk new_AGEMA_reg_buffer_7729 ( .C (clk), .D (new_AGEMA_signal_20452), .Q (new_AGEMA_signal_20453) ) ;
    buf_clk new_AGEMA_reg_buffer_7732 ( .C (clk), .D (new_AGEMA_signal_20455), .Q (new_AGEMA_signal_20456) ) ;
    buf_clk new_AGEMA_reg_buffer_7735 ( .C (clk), .D (new_AGEMA_signal_20458), .Q (new_AGEMA_signal_20459) ) ;
    buf_clk new_AGEMA_reg_buffer_7738 ( .C (clk), .D (new_AGEMA_signal_20461), .Q (new_AGEMA_signal_20462) ) ;
    buf_clk new_AGEMA_reg_buffer_7741 ( .C (clk), .D (new_AGEMA_signal_20464), .Q (new_AGEMA_signal_20465) ) ;
    buf_clk new_AGEMA_reg_buffer_7744 ( .C (clk), .D (new_AGEMA_signal_20467), .Q (new_AGEMA_signal_20468) ) ;
    buf_clk new_AGEMA_reg_buffer_7747 ( .C (clk), .D (new_AGEMA_signal_20470), .Q (new_AGEMA_signal_20471) ) ;
    buf_clk new_AGEMA_reg_buffer_7750 ( .C (clk), .D (new_AGEMA_signal_20473), .Q (new_AGEMA_signal_20474) ) ;
    buf_clk new_AGEMA_reg_buffer_7753 ( .C (clk), .D (new_AGEMA_signal_20476), .Q (new_AGEMA_signal_20477) ) ;
    buf_clk new_AGEMA_reg_buffer_7756 ( .C (clk), .D (new_AGEMA_signal_20479), .Q (new_AGEMA_signal_20480) ) ;
    buf_clk new_AGEMA_reg_buffer_7759 ( .C (clk), .D (new_AGEMA_signal_20482), .Q (new_AGEMA_signal_20483) ) ;
    buf_clk new_AGEMA_reg_buffer_7762 ( .C (clk), .D (new_AGEMA_signal_20485), .Q (new_AGEMA_signal_20486) ) ;
    buf_clk new_AGEMA_reg_buffer_7765 ( .C (clk), .D (new_AGEMA_signal_20488), .Q (new_AGEMA_signal_20489) ) ;
    buf_clk new_AGEMA_reg_buffer_7768 ( .C (clk), .D (new_AGEMA_signal_20491), .Q (new_AGEMA_signal_20492) ) ;
    buf_clk new_AGEMA_reg_buffer_7771 ( .C (clk), .D (new_AGEMA_signal_20494), .Q (new_AGEMA_signal_20495) ) ;
    buf_clk new_AGEMA_reg_buffer_7774 ( .C (clk), .D (new_AGEMA_signal_20497), .Q (new_AGEMA_signal_20498) ) ;
    buf_clk new_AGEMA_reg_buffer_7777 ( .C (clk), .D (new_AGEMA_signal_20500), .Q (new_AGEMA_signal_20501) ) ;
    buf_clk new_AGEMA_reg_buffer_7780 ( .C (clk), .D (new_AGEMA_signal_20503), .Q (new_AGEMA_signal_20504) ) ;
    buf_clk new_AGEMA_reg_buffer_7783 ( .C (clk), .D (new_AGEMA_signal_20506), .Q (new_AGEMA_signal_20507) ) ;
    buf_clk new_AGEMA_reg_buffer_7786 ( .C (clk), .D (new_AGEMA_signal_20509), .Q (new_AGEMA_signal_20510) ) ;
    buf_clk new_AGEMA_reg_buffer_7789 ( .C (clk), .D (new_AGEMA_signal_20512), .Q (new_AGEMA_signal_20513) ) ;
    buf_clk new_AGEMA_reg_buffer_7792 ( .C (clk), .D (new_AGEMA_signal_20515), .Q (new_AGEMA_signal_20516) ) ;
    buf_clk new_AGEMA_reg_buffer_7795 ( .C (clk), .D (new_AGEMA_signal_20518), .Q (new_AGEMA_signal_20519) ) ;
    buf_clk new_AGEMA_reg_buffer_7798 ( .C (clk), .D (new_AGEMA_signal_20521), .Q (new_AGEMA_signal_20522) ) ;
    buf_clk new_AGEMA_reg_buffer_7801 ( .C (clk), .D (new_AGEMA_signal_20524), .Q (new_AGEMA_signal_20525) ) ;
    buf_clk new_AGEMA_reg_buffer_7804 ( .C (clk), .D (new_AGEMA_signal_20527), .Q (new_AGEMA_signal_20528) ) ;
    buf_clk new_AGEMA_reg_buffer_7807 ( .C (clk), .D (new_AGEMA_signal_20530), .Q (new_AGEMA_signal_20531) ) ;
    buf_clk new_AGEMA_reg_buffer_7810 ( .C (clk), .D (new_AGEMA_signal_20533), .Q (new_AGEMA_signal_20534) ) ;
    buf_clk new_AGEMA_reg_buffer_7813 ( .C (clk), .D (new_AGEMA_signal_20536), .Q (new_AGEMA_signal_20537) ) ;
    buf_clk new_AGEMA_reg_buffer_7816 ( .C (clk), .D (new_AGEMA_signal_20539), .Q (new_AGEMA_signal_20540) ) ;
    buf_clk new_AGEMA_reg_buffer_7819 ( .C (clk), .D (new_AGEMA_signal_20542), .Q (new_AGEMA_signal_20543) ) ;
    buf_clk new_AGEMA_reg_buffer_7822 ( .C (clk), .D (new_AGEMA_signal_20545), .Q (new_AGEMA_signal_20546) ) ;
    buf_clk new_AGEMA_reg_buffer_7825 ( .C (clk), .D (new_AGEMA_signal_20548), .Q (new_AGEMA_signal_20549) ) ;
    buf_clk new_AGEMA_reg_buffer_7828 ( .C (clk), .D (new_AGEMA_signal_20551), .Q (new_AGEMA_signal_20552) ) ;
    buf_clk new_AGEMA_reg_buffer_7831 ( .C (clk), .D (new_AGEMA_signal_20554), .Q (new_AGEMA_signal_20555) ) ;
    buf_clk new_AGEMA_reg_buffer_7834 ( .C (clk), .D (new_AGEMA_signal_20557), .Q (new_AGEMA_signal_20558) ) ;
    buf_clk new_AGEMA_reg_buffer_7837 ( .C (clk), .D (new_AGEMA_signal_20560), .Q (new_AGEMA_signal_20561) ) ;
    buf_clk new_AGEMA_reg_buffer_7840 ( .C (clk), .D (new_AGEMA_signal_20563), .Q (new_AGEMA_signal_20564) ) ;
    buf_clk new_AGEMA_reg_buffer_7843 ( .C (clk), .D (new_AGEMA_signal_20566), .Q (new_AGEMA_signal_20567) ) ;
    buf_clk new_AGEMA_reg_buffer_7846 ( .C (clk), .D (new_AGEMA_signal_20569), .Q (new_AGEMA_signal_20570) ) ;
    buf_clk new_AGEMA_reg_buffer_7849 ( .C (clk), .D (new_AGEMA_signal_20572), .Q (new_AGEMA_signal_20573) ) ;
    buf_clk new_AGEMA_reg_buffer_7852 ( .C (clk), .D (new_AGEMA_signal_20575), .Q (new_AGEMA_signal_20576) ) ;
    buf_clk new_AGEMA_reg_buffer_7855 ( .C (clk), .D (new_AGEMA_signal_20578), .Q (new_AGEMA_signal_20579) ) ;
    buf_clk new_AGEMA_reg_buffer_7858 ( .C (clk), .D (new_AGEMA_signal_20581), .Q (new_AGEMA_signal_20582) ) ;
    buf_clk new_AGEMA_reg_buffer_7861 ( .C (clk), .D (new_AGEMA_signal_20584), .Q (new_AGEMA_signal_20585) ) ;
    buf_clk new_AGEMA_reg_buffer_7864 ( .C (clk), .D (new_AGEMA_signal_20587), .Q (new_AGEMA_signal_20588) ) ;
    buf_clk new_AGEMA_reg_buffer_7867 ( .C (clk), .D (new_AGEMA_signal_20590), .Q (new_AGEMA_signal_20591) ) ;
    buf_clk new_AGEMA_reg_buffer_7870 ( .C (clk), .D (new_AGEMA_signal_20593), .Q (new_AGEMA_signal_20594) ) ;
    buf_clk new_AGEMA_reg_buffer_7873 ( .C (clk), .D (new_AGEMA_signal_20596), .Q (new_AGEMA_signal_20597) ) ;
    buf_clk new_AGEMA_reg_buffer_7876 ( .C (clk), .D (new_AGEMA_signal_20599), .Q (new_AGEMA_signal_20600) ) ;
    buf_clk new_AGEMA_reg_buffer_7879 ( .C (clk), .D (new_AGEMA_signal_20602), .Q (new_AGEMA_signal_20603) ) ;
    buf_clk new_AGEMA_reg_buffer_7882 ( .C (clk), .D (new_AGEMA_signal_20605), .Q (new_AGEMA_signal_20606) ) ;
    buf_clk new_AGEMA_reg_buffer_7885 ( .C (clk), .D (new_AGEMA_signal_20608), .Q (new_AGEMA_signal_20609) ) ;
    buf_clk new_AGEMA_reg_buffer_7888 ( .C (clk), .D (new_AGEMA_signal_20611), .Q (new_AGEMA_signal_20612) ) ;
    buf_clk new_AGEMA_reg_buffer_7891 ( .C (clk), .D (new_AGEMA_signal_20614), .Q (new_AGEMA_signal_20615) ) ;
    buf_clk new_AGEMA_reg_buffer_7894 ( .C (clk), .D (new_AGEMA_signal_20617), .Q (new_AGEMA_signal_20618) ) ;
    buf_clk new_AGEMA_reg_buffer_7897 ( .C (clk), .D (new_AGEMA_signal_20620), .Q (new_AGEMA_signal_20621) ) ;
    buf_clk new_AGEMA_reg_buffer_7900 ( .C (clk), .D (new_AGEMA_signal_20623), .Q (new_AGEMA_signal_20624) ) ;
    buf_clk new_AGEMA_reg_buffer_7903 ( .C (clk), .D (new_AGEMA_signal_20626), .Q (new_AGEMA_signal_20627) ) ;
    buf_clk new_AGEMA_reg_buffer_7906 ( .C (clk), .D (new_AGEMA_signal_20629), .Q (new_AGEMA_signal_20630) ) ;
    buf_clk new_AGEMA_reg_buffer_7909 ( .C (clk), .D (new_AGEMA_signal_20632), .Q (new_AGEMA_signal_20633) ) ;
    buf_clk new_AGEMA_reg_buffer_7912 ( .C (clk), .D (new_AGEMA_signal_20635), .Q (new_AGEMA_signal_20636) ) ;
    buf_clk new_AGEMA_reg_buffer_7915 ( .C (clk), .D (new_AGEMA_signal_20638), .Q (new_AGEMA_signal_20639) ) ;
    buf_clk new_AGEMA_reg_buffer_7918 ( .C (clk), .D (new_AGEMA_signal_20641), .Q (new_AGEMA_signal_20642) ) ;
    buf_clk new_AGEMA_reg_buffer_7921 ( .C (clk), .D (new_AGEMA_signal_20644), .Q (new_AGEMA_signal_20645) ) ;
    buf_clk new_AGEMA_reg_buffer_7924 ( .C (clk), .D (new_AGEMA_signal_20647), .Q (new_AGEMA_signal_20648) ) ;
    buf_clk new_AGEMA_reg_buffer_7927 ( .C (clk), .D (new_AGEMA_signal_20650), .Q (new_AGEMA_signal_20651) ) ;
    buf_clk new_AGEMA_reg_buffer_7930 ( .C (clk), .D (new_AGEMA_signal_20653), .Q (new_AGEMA_signal_20654) ) ;
    buf_clk new_AGEMA_reg_buffer_7933 ( .C (clk), .D (new_AGEMA_signal_20656), .Q (new_AGEMA_signal_20657) ) ;
    buf_clk new_AGEMA_reg_buffer_7936 ( .C (clk), .D (new_AGEMA_signal_20659), .Q (new_AGEMA_signal_20660) ) ;
    buf_clk new_AGEMA_reg_buffer_7939 ( .C (clk), .D (new_AGEMA_signal_20662), .Q (new_AGEMA_signal_20663) ) ;
    buf_clk new_AGEMA_reg_buffer_7942 ( .C (clk), .D (new_AGEMA_signal_20665), .Q (new_AGEMA_signal_20666) ) ;
    buf_clk new_AGEMA_reg_buffer_7945 ( .C (clk), .D (new_AGEMA_signal_20668), .Q (new_AGEMA_signal_20669) ) ;
    buf_clk new_AGEMA_reg_buffer_7948 ( .C (clk), .D (new_AGEMA_signal_20671), .Q (new_AGEMA_signal_20672) ) ;
    buf_clk new_AGEMA_reg_buffer_7951 ( .C (clk), .D (new_AGEMA_signal_20674), .Q (new_AGEMA_signal_20675) ) ;
    buf_clk new_AGEMA_reg_buffer_7954 ( .C (clk), .D (new_AGEMA_signal_20677), .Q (new_AGEMA_signal_20678) ) ;
    buf_clk new_AGEMA_reg_buffer_7957 ( .C (clk), .D (new_AGEMA_signal_20680), .Q (new_AGEMA_signal_20681) ) ;
    buf_clk new_AGEMA_reg_buffer_7960 ( .C (clk), .D (new_AGEMA_signal_20683), .Q (new_AGEMA_signal_20684) ) ;
    buf_clk new_AGEMA_reg_buffer_7963 ( .C (clk), .D (new_AGEMA_signal_20686), .Q (new_AGEMA_signal_20687) ) ;
    buf_clk new_AGEMA_reg_buffer_7966 ( .C (clk), .D (new_AGEMA_signal_20689), .Q (new_AGEMA_signal_20690) ) ;
    buf_clk new_AGEMA_reg_buffer_7969 ( .C (clk), .D (new_AGEMA_signal_20692), .Q (new_AGEMA_signal_20693) ) ;
    buf_clk new_AGEMA_reg_buffer_7972 ( .C (clk), .D (new_AGEMA_signal_20695), .Q (new_AGEMA_signal_20696) ) ;
    buf_clk new_AGEMA_reg_buffer_7975 ( .C (clk), .D (new_AGEMA_signal_20698), .Q (new_AGEMA_signal_20699) ) ;
    buf_clk new_AGEMA_reg_buffer_7978 ( .C (clk), .D (new_AGEMA_signal_20701), .Q (new_AGEMA_signal_20702) ) ;
    buf_clk new_AGEMA_reg_buffer_7981 ( .C (clk), .D (new_AGEMA_signal_20704), .Q (new_AGEMA_signal_20705) ) ;
    buf_clk new_AGEMA_reg_buffer_7984 ( .C (clk), .D (new_AGEMA_signal_20707), .Q (new_AGEMA_signal_20708) ) ;
    buf_clk new_AGEMA_reg_buffer_7987 ( .C (clk), .D (new_AGEMA_signal_20710), .Q (new_AGEMA_signal_20711) ) ;
    buf_clk new_AGEMA_reg_buffer_7990 ( .C (clk), .D (new_AGEMA_signal_20713), .Q (new_AGEMA_signal_20714) ) ;
    buf_clk new_AGEMA_reg_buffer_7993 ( .C (clk), .D (new_AGEMA_signal_20716), .Q (new_AGEMA_signal_20717) ) ;
    buf_clk new_AGEMA_reg_buffer_7996 ( .C (clk), .D (new_AGEMA_signal_20719), .Q (new_AGEMA_signal_20720) ) ;
    buf_clk new_AGEMA_reg_buffer_7999 ( .C (clk), .D (new_AGEMA_signal_20722), .Q (new_AGEMA_signal_20723) ) ;
    buf_clk new_AGEMA_reg_buffer_8002 ( .C (clk), .D (new_AGEMA_signal_20725), .Q (new_AGEMA_signal_20726) ) ;
    buf_clk new_AGEMA_reg_buffer_8005 ( .C (clk), .D (new_AGEMA_signal_20728), .Q (new_AGEMA_signal_20729) ) ;
    buf_clk new_AGEMA_reg_buffer_8008 ( .C (clk), .D (new_AGEMA_signal_20731), .Q (new_AGEMA_signal_20732) ) ;
    buf_clk new_AGEMA_reg_buffer_8011 ( .C (clk), .D (new_AGEMA_signal_20734), .Q (new_AGEMA_signal_20735) ) ;
    buf_clk new_AGEMA_reg_buffer_8014 ( .C (clk), .D (new_AGEMA_signal_20737), .Q (new_AGEMA_signal_20738) ) ;
    buf_clk new_AGEMA_reg_buffer_8017 ( .C (clk), .D (new_AGEMA_signal_20740), .Q (new_AGEMA_signal_20741) ) ;
    buf_clk new_AGEMA_reg_buffer_8020 ( .C (clk), .D (new_AGEMA_signal_20743), .Q (new_AGEMA_signal_20744) ) ;
    buf_clk new_AGEMA_reg_buffer_8023 ( .C (clk), .D (new_AGEMA_signal_20746), .Q (new_AGEMA_signal_20747) ) ;
    buf_clk new_AGEMA_reg_buffer_8026 ( .C (clk), .D (new_AGEMA_signal_20749), .Q (new_AGEMA_signal_20750) ) ;
    buf_clk new_AGEMA_reg_buffer_8029 ( .C (clk), .D (new_AGEMA_signal_20752), .Q (new_AGEMA_signal_20753) ) ;
    buf_clk new_AGEMA_reg_buffer_8032 ( .C (clk), .D (new_AGEMA_signal_20755), .Q (new_AGEMA_signal_20756) ) ;
    buf_clk new_AGEMA_reg_buffer_8035 ( .C (clk), .D (new_AGEMA_signal_20758), .Q (new_AGEMA_signal_20759) ) ;
    buf_clk new_AGEMA_reg_buffer_8038 ( .C (clk), .D (new_AGEMA_signal_20761), .Q (new_AGEMA_signal_20762) ) ;
    buf_clk new_AGEMA_reg_buffer_8041 ( .C (clk), .D (new_AGEMA_signal_20764), .Q (new_AGEMA_signal_20765) ) ;
    buf_clk new_AGEMA_reg_buffer_8044 ( .C (clk), .D (new_AGEMA_signal_20767), .Q (new_AGEMA_signal_20768) ) ;
    buf_clk new_AGEMA_reg_buffer_8047 ( .C (clk), .D (new_AGEMA_signal_20770), .Q (new_AGEMA_signal_20771) ) ;
    buf_clk new_AGEMA_reg_buffer_8050 ( .C (clk), .D (new_AGEMA_signal_20773), .Q (new_AGEMA_signal_20774) ) ;
    buf_clk new_AGEMA_reg_buffer_8053 ( .C (clk), .D (new_AGEMA_signal_20776), .Q (new_AGEMA_signal_20777) ) ;
    buf_clk new_AGEMA_reg_buffer_8056 ( .C (clk), .D (new_AGEMA_signal_20779), .Q (new_AGEMA_signal_20780) ) ;
    buf_clk new_AGEMA_reg_buffer_8059 ( .C (clk), .D (new_AGEMA_signal_20782), .Q (new_AGEMA_signal_20783) ) ;
    buf_clk new_AGEMA_reg_buffer_8062 ( .C (clk), .D (new_AGEMA_signal_20785), .Q (new_AGEMA_signal_20786) ) ;
    buf_clk new_AGEMA_reg_buffer_8065 ( .C (clk), .D (new_AGEMA_signal_20788), .Q (new_AGEMA_signal_20789) ) ;
    buf_clk new_AGEMA_reg_buffer_8068 ( .C (clk), .D (new_AGEMA_signal_20791), .Q (new_AGEMA_signal_20792) ) ;
    buf_clk new_AGEMA_reg_buffer_8071 ( .C (clk), .D (new_AGEMA_signal_20794), .Q (new_AGEMA_signal_20795) ) ;
    buf_clk new_AGEMA_reg_buffer_8074 ( .C (clk), .D (new_AGEMA_signal_20797), .Q (new_AGEMA_signal_20798) ) ;
    buf_clk new_AGEMA_reg_buffer_8077 ( .C (clk), .D (new_AGEMA_signal_20800), .Q (new_AGEMA_signal_20801) ) ;
    buf_clk new_AGEMA_reg_buffer_8080 ( .C (clk), .D (new_AGEMA_signal_20803), .Q (new_AGEMA_signal_20804) ) ;
    buf_clk new_AGEMA_reg_buffer_8083 ( .C (clk), .D (new_AGEMA_signal_20806), .Q (new_AGEMA_signal_20807) ) ;
    buf_clk new_AGEMA_reg_buffer_8086 ( .C (clk), .D (new_AGEMA_signal_20809), .Q (new_AGEMA_signal_20810) ) ;
    buf_clk new_AGEMA_reg_buffer_8089 ( .C (clk), .D (new_AGEMA_signal_20812), .Q (new_AGEMA_signal_20813) ) ;
    buf_clk new_AGEMA_reg_buffer_8092 ( .C (clk), .D (new_AGEMA_signal_20815), .Q (new_AGEMA_signal_20816) ) ;
    buf_clk new_AGEMA_reg_buffer_8095 ( .C (clk), .D (new_AGEMA_signal_20818), .Q (new_AGEMA_signal_20819) ) ;
    buf_clk new_AGEMA_reg_buffer_8098 ( .C (clk), .D (new_AGEMA_signal_20821), .Q (new_AGEMA_signal_20822) ) ;
    buf_clk new_AGEMA_reg_buffer_8101 ( .C (clk), .D (new_AGEMA_signal_20824), .Q (new_AGEMA_signal_20825) ) ;
    buf_clk new_AGEMA_reg_buffer_8104 ( .C (clk), .D (new_AGEMA_signal_20827), .Q (new_AGEMA_signal_20828) ) ;
    buf_clk new_AGEMA_reg_buffer_8107 ( .C (clk), .D (new_AGEMA_signal_20830), .Q (new_AGEMA_signal_20831) ) ;
    buf_clk new_AGEMA_reg_buffer_8110 ( .C (clk), .D (new_AGEMA_signal_20833), .Q (new_AGEMA_signal_20834) ) ;
    buf_clk new_AGEMA_reg_buffer_8113 ( .C (clk), .D (new_AGEMA_signal_20836), .Q (new_AGEMA_signal_20837) ) ;
    buf_clk new_AGEMA_reg_buffer_8116 ( .C (clk), .D (new_AGEMA_signal_20839), .Q (new_AGEMA_signal_20840) ) ;
    buf_clk new_AGEMA_reg_buffer_8119 ( .C (clk), .D (new_AGEMA_signal_20842), .Q (new_AGEMA_signal_20843) ) ;
    buf_clk new_AGEMA_reg_buffer_8122 ( .C (clk), .D (new_AGEMA_signal_20845), .Q (new_AGEMA_signal_20846) ) ;
    buf_clk new_AGEMA_reg_buffer_8125 ( .C (clk), .D (new_AGEMA_signal_20848), .Q (new_AGEMA_signal_20849) ) ;
    buf_clk new_AGEMA_reg_buffer_8128 ( .C (clk), .D (new_AGEMA_signal_20851), .Q (new_AGEMA_signal_20852) ) ;
    buf_clk new_AGEMA_reg_buffer_8131 ( .C (clk), .D (new_AGEMA_signal_20854), .Q (new_AGEMA_signal_20855) ) ;
    buf_clk new_AGEMA_reg_buffer_8134 ( .C (clk), .D (new_AGEMA_signal_20857), .Q (new_AGEMA_signal_20858) ) ;
    buf_clk new_AGEMA_reg_buffer_8137 ( .C (clk), .D (new_AGEMA_signal_20860), .Q (new_AGEMA_signal_20861) ) ;
    buf_clk new_AGEMA_reg_buffer_8140 ( .C (clk), .D (new_AGEMA_signal_20863), .Q (new_AGEMA_signal_20864) ) ;
    buf_clk new_AGEMA_reg_buffer_8143 ( .C (clk), .D (new_AGEMA_signal_20866), .Q (new_AGEMA_signal_20867) ) ;
    buf_clk new_AGEMA_reg_buffer_8146 ( .C (clk), .D (new_AGEMA_signal_20869), .Q (new_AGEMA_signal_20870) ) ;
    buf_clk new_AGEMA_reg_buffer_8149 ( .C (clk), .D (new_AGEMA_signal_20872), .Q (new_AGEMA_signal_20873) ) ;
    buf_clk new_AGEMA_reg_buffer_8152 ( .C (clk), .D (new_AGEMA_signal_20875), .Q (new_AGEMA_signal_20876) ) ;
    buf_clk new_AGEMA_reg_buffer_8155 ( .C (clk), .D (new_AGEMA_signal_20878), .Q (new_AGEMA_signal_20879) ) ;
    buf_clk new_AGEMA_reg_buffer_8158 ( .C (clk), .D (new_AGEMA_signal_20881), .Q (new_AGEMA_signal_20882) ) ;
    buf_clk new_AGEMA_reg_buffer_8161 ( .C (clk), .D (new_AGEMA_signal_20884), .Q (new_AGEMA_signal_20885) ) ;
    buf_clk new_AGEMA_reg_buffer_8164 ( .C (clk), .D (new_AGEMA_signal_20887), .Q (new_AGEMA_signal_20888) ) ;
    buf_clk new_AGEMA_reg_buffer_8167 ( .C (clk), .D (new_AGEMA_signal_20890), .Q (new_AGEMA_signal_20891) ) ;
    buf_clk new_AGEMA_reg_buffer_8170 ( .C (clk), .D (new_AGEMA_signal_20893), .Q (new_AGEMA_signal_20894) ) ;
    buf_clk new_AGEMA_reg_buffer_8173 ( .C (clk), .D (new_AGEMA_signal_20896), .Q (new_AGEMA_signal_20897) ) ;
    buf_clk new_AGEMA_reg_buffer_8176 ( .C (clk), .D (new_AGEMA_signal_20899), .Q (new_AGEMA_signal_20900) ) ;
    buf_clk new_AGEMA_reg_buffer_8179 ( .C (clk), .D (new_AGEMA_signal_20902), .Q (new_AGEMA_signal_20903) ) ;
    buf_clk new_AGEMA_reg_buffer_8182 ( .C (clk), .D (new_AGEMA_signal_20905), .Q (new_AGEMA_signal_20906) ) ;
    buf_clk new_AGEMA_reg_buffer_8185 ( .C (clk), .D (new_AGEMA_signal_20908), .Q (new_AGEMA_signal_20909) ) ;
    buf_clk new_AGEMA_reg_buffer_8188 ( .C (clk), .D (new_AGEMA_signal_20911), .Q (new_AGEMA_signal_20912) ) ;
    buf_clk new_AGEMA_reg_buffer_8191 ( .C (clk), .D (new_AGEMA_signal_20914), .Q (new_AGEMA_signal_20915) ) ;
    buf_clk new_AGEMA_reg_buffer_8194 ( .C (clk), .D (new_AGEMA_signal_20917), .Q (new_AGEMA_signal_20918) ) ;
    buf_clk new_AGEMA_reg_buffer_8197 ( .C (clk), .D (new_AGEMA_signal_20920), .Q (new_AGEMA_signal_20921) ) ;
    buf_clk new_AGEMA_reg_buffer_8200 ( .C (clk), .D (new_AGEMA_signal_20923), .Q (new_AGEMA_signal_20924) ) ;
    buf_clk new_AGEMA_reg_buffer_8203 ( .C (clk), .D (new_AGEMA_signal_20926), .Q (new_AGEMA_signal_20927) ) ;
    buf_clk new_AGEMA_reg_buffer_8206 ( .C (clk), .D (new_AGEMA_signal_20929), .Q (new_AGEMA_signal_20930) ) ;
    buf_clk new_AGEMA_reg_buffer_8209 ( .C (clk), .D (new_AGEMA_signal_20932), .Q (new_AGEMA_signal_20933) ) ;
    buf_clk new_AGEMA_reg_buffer_8212 ( .C (clk), .D (new_AGEMA_signal_20935), .Q (new_AGEMA_signal_20936) ) ;
    buf_clk new_AGEMA_reg_buffer_8215 ( .C (clk), .D (new_AGEMA_signal_20938), .Q (new_AGEMA_signal_20939) ) ;
    buf_clk new_AGEMA_reg_buffer_8218 ( .C (clk), .D (new_AGEMA_signal_20941), .Q (new_AGEMA_signal_20942) ) ;
    buf_clk new_AGEMA_reg_buffer_8221 ( .C (clk), .D (new_AGEMA_signal_20944), .Q (new_AGEMA_signal_20945) ) ;
    buf_clk new_AGEMA_reg_buffer_8224 ( .C (clk), .D (new_AGEMA_signal_20947), .Q (new_AGEMA_signal_20948) ) ;
    buf_clk new_AGEMA_reg_buffer_8227 ( .C (clk), .D (new_AGEMA_signal_20950), .Q (new_AGEMA_signal_20951) ) ;
    buf_clk new_AGEMA_reg_buffer_8230 ( .C (clk), .D (new_AGEMA_signal_20953), .Q (new_AGEMA_signal_20954) ) ;
    buf_clk new_AGEMA_reg_buffer_8233 ( .C (clk), .D (new_AGEMA_signal_20956), .Q (new_AGEMA_signal_20957) ) ;
    buf_clk new_AGEMA_reg_buffer_8236 ( .C (clk), .D (new_AGEMA_signal_20959), .Q (new_AGEMA_signal_20960) ) ;
    buf_clk new_AGEMA_reg_buffer_8239 ( .C (clk), .D (new_AGEMA_signal_20962), .Q (new_AGEMA_signal_20963) ) ;
    buf_clk new_AGEMA_reg_buffer_8242 ( .C (clk), .D (new_AGEMA_signal_20965), .Q (new_AGEMA_signal_20966) ) ;
    buf_clk new_AGEMA_reg_buffer_8245 ( .C (clk), .D (new_AGEMA_signal_20968), .Q (new_AGEMA_signal_20969) ) ;
    buf_clk new_AGEMA_reg_buffer_8248 ( .C (clk), .D (new_AGEMA_signal_20971), .Q (new_AGEMA_signal_20972) ) ;
    buf_clk new_AGEMA_reg_buffer_8251 ( .C (clk), .D (new_AGEMA_signal_20974), .Q (new_AGEMA_signal_20975) ) ;
    buf_clk new_AGEMA_reg_buffer_8254 ( .C (clk), .D (new_AGEMA_signal_20977), .Q (new_AGEMA_signal_20978) ) ;
    buf_clk new_AGEMA_reg_buffer_8257 ( .C (clk), .D (new_AGEMA_signal_20980), .Q (new_AGEMA_signal_20981) ) ;
    buf_clk new_AGEMA_reg_buffer_8260 ( .C (clk), .D (new_AGEMA_signal_20983), .Q (new_AGEMA_signal_20984) ) ;
    buf_clk new_AGEMA_reg_buffer_8263 ( .C (clk), .D (new_AGEMA_signal_20986), .Q (new_AGEMA_signal_20987) ) ;
    buf_clk new_AGEMA_reg_buffer_8266 ( .C (clk), .D (new_AGEMA_signal_20989), .Q (new_AGEMA_signal_20990) ) ;
    buf_clk new_AGEMA_reg_buffer_8269 ( .C (clk), .D (new_AGEMA_signal_20992), .Q (new_AGEMA_signal_20993) ) ;
    buf_clk new_AGEMA_reg_buffer_8272 ( .C (clk), .D (new_AGEMA_signal_20995), .Q (new_AGEMA_signal_20996) ) ;
    buf_clk new_AGEMA_reg_buffer_8275 ( .C (clk), .D (new_AGEMA_signal_20998), .Q (new_AGEMA_signal_20999) ) ;
    buf_clk new_AGEMA_reg_buffer_8278 ( .C (clk), .D (new_AGEMA_signal_21001), .Q (new_AGEMA_signal_21002) ) ;
    buf_clk new_AGEMA_reg_buffer_8281 ( .C (clk), .D (new_AGEMA_signal_21004), .Q (new_AGEMA_signal_21005) ) ;
    buf_clk new_AGEMA_reg_buffer_8284 ( .C (clk), .D (new_AGEMA_signal_21007), .Q (new_AGEMA_signal_21008) ) ;
    buf_clk new_AGEMA_reg_buffer_8287 ( .C (clk), .D (new_AGEMA_signal_21010), .Q (new_AGEMA_signal_21011) ) ;
    buf_clk new_AGEMA_reg_buffer_8290 ( .C (clk), .D (new_AGEMA_signal_21013), .Q (new_AGEMA_signal_21014) ) ;
    buf_clk new_AGEMA_reg_buffer_8293 ( .C (clk), .D (new_AGEMA_signal_21016), .Q (new_AGEMA_signal_21017) ) ;
    buf_clk new_AGEMA_reg_buffer_8296 ( .C (clk), .D (new_AGEMA_signal_21019), .Q (new_AGEMA_signal_21020) ) ;
    buf_clk new_AGEMA_reg_buffer_8299 ( .C (clk), .D (new_AGEMA_signal_21022), .Q (new_AGEMA_signal_21023) ) ;
    buf_clk new_AGEMA_reg_buffer_8302 ( .C (clk), .D (new_AGEMA_signal_21025), .Q (new_AGEMA_signal_21026) ) ;
    buf_clk new_AGEMA_reg_buffer_8305 ( .C (clk), .D (new_AGEMA_signal_21028), .Q (new_AGEMA_signal_21029) ) ;
    buf_clk new_AGEMA_reg_buffer_8308 ( .C (clk), .D (new_AGEMA_signal_21031), .Q (new_AGEMA_signal_21032) ) ;
    buf_clk new_AGEMA_reg_buffer_8311 ( .C (clk), .D (new_AGEMA_signal_21034), .Q (new_AGEMA_signal_21035) ) ;
    buf_clk new_AGEMA_reg_buffer_8314 ( .C (clk), .D (new_AGEMA_signal_21037), .Q (new_AGEMA_signal_21038) ) ;
    buf_clk new_AGEMA_reg_buffer_8317 ( .C (clk), .D (new_AGEMA_signal_21040), .Q (new_AGEMA_signal_21041) ) ;
    buf_clk new_AGEMA_reg_buffer_8320 ( .C (clk), .D (new_AGEMA_signal_21043), .Q (new_AGEMA_signal_21044) ) ;
    buf_clk new_AGEMA_reg_buffer_8323 ( .C (clk), .D (new_AGEMA_signal_21046), .Q (new_AGEMA_signal_21047) ) ;
    buf_clk new_AGEMA_reg_buffer_8326 ( .C (clk), .D (new_AGEMA_signal_21049), .Q (new_AGEMA_signal_21050) ) ;
    buf_clk new_AGEMA_reg_buffer_8329 ( .C (clk), .D (new_AGEMA_signal_21052), .Q (new_AGEMA_signal_21053) ) ;
    buf_clk new_AGEMA_reg_buffer_8332 ( .C (clk), .D (new_AGEMA_signal_21055), .Q (new_AGEMA_signal_21056) ) ;
    buf_clk new_AGEMA_reg_buffer_8335 ( .C (clk), .D (new_AGEMA_signal_21058), .Q (new_AGEMA_signal_21059) ) ;
    buf_clk new_AGEMA_reg_buffer_8338 ( .C (clk), .D (new_AGEMA_signal_21061), .Q (new_AGEMA_signal_21062) ) ;
    buf_clk new_AGEMA_reg_buffer_8341 ( .C (clk), .D (new_AGEMA_signal_21064), .Q (new_AGEMA_signal_21065) ) ;
    buf_clk new_AGEMA_reg_buffer_8344 ( .C (clk), .D (new_AGEMA_signal_21067), .Q (new_AGEMA_signal_21068) ) ;
    buf_clk new_AGEMA_reg_buffer_8347 ( .C (clk), .D (new_AGEMA_signal_21070), .Q (new_AGEMA_signal_21071) ) ;
    buf_clk new_AGEMA_reg_buffer_8350 ( .C (clk), .D (new_AGEMA_signal_21073), .Q (new_AGEMA_signal_21074) ) ;
    buf_clk new_AGEMA_reg_buffer_8353 ( .C (clk), .D (new_AGEMA_signal_21076), .Q (new_AGEMA_signal_21077) ) ;
    buf_clk new_AGEMA_reg_buffer_8356 ( .C (clk), .D (new_AGEMA_signal_21079), .Q (new_AGEMA_signal_21080) ) ;
    buf_clk new_AGEMA_reg_buffer_8359 ( .C (clk), .D (new_AGEMA_signal_21082), .Q (new_AGEMA_signal_21083) ) ;
    buf_clk new_AGEMA_reg_buffer_8362 ( .C (clk), .D (new_AGEMA_signal_21085), .Q (new_AGEMA_signal_21086) ) ;
    buf_clk new_AGEMA_reg_buffer_8365 ( .C (clk), .D (new_AGEMA_signal_21088), .Q (new_AGEMA_signal_21089) ) ;
    buf_clk new_AGEMA_reg_buffer_8368 ( .C (clk), .D (new_AGEMA_signal_21091), .Q (new_AGEMA_signal_21092) ) ;
    buf_clk new_AGEMA_reg_buffer_8371 ( .C (clk), .D (new_AGEMA_signal_21094), .Q (new_AGEMA_signal_21095) ) ;
    buf_clk new_AGEMA_reg_buffer_8374 ( .C (clk), .D (new_AGEMA_signal_21097), .Q (new_AGEMA_signal_21098) ) ;
    buf_clk new_AGEMA_reg_buffer_8377 ( .C (clk), .D (new_AGEMA_signal_21100), .Q (new_AGEMA_signal_21101) ) ;
    buf_clk new_AGEMA_reg_buffer_8380 ( .C (clk), .D (new_AGEMA_signal_21103), .Q (new_AGEMA_signal_21104) ) ;
    buf_clk new_AGEMA_reg_buffer_8383 ( .C (clk), .D (new_AGEMA_signal_21106), .Q (new_AGEMA_signal_21107) ) ;
    buf_clk new_AGEMA_reg_buffer_8386 ( .C (clk), .D (new_AGEMA_signal_21109), .Q (new_AGEMA_signal_21110) ) ;
    buf_clk new_AGEMA_reg_buffer_8389 ( .C (clk), .D (new_AGEMA_signal_21112), .Q (new_AGEMA_signal_21113) ) ;
    buf_clk new_AGEMA_reg_buffer_8392 ( .C (clk), .D (new_AGEMA_signal_21115), .Q (new_AGEMA_signal_21116) ) ;
    buf_clk new_AGEMA_reg_buffer_8395 ( .C (clk), .D (new_AGEMA_signal_21118), .Q (new_AGEMA_signal_21119) ) ;
    buf_clk new_AGEMA_reg_buffer_8398 ( .C (clk), .D (new_AGEMA_signal_21121), .Q (new_AGEMA_signal_21122) ) ;
    buf_clk new_AGEMA_reg_buffer_8401 ( .C (clk), .D (new_AGEMA_signal_21124), .Q (new_AGEMA_signal_21125) ) ;
    buf_clk new_AGEMA_reg_buffer_8404 ( .C (clk), .D (new_AGEMA_signal_21127), .Q (new_AGEMA_signal_21128) ) ;
    buf_clk new_AGEMA_reg_buffer_8407 ( .C (clk), .D (new_AGEMA_signal_21130), .Q (new_AGEMA_signal_21131) ) ;
    buf_clk new_AGEMA_reg_buffer_8410 ( .C (clk), .D (new_AGEMA_signal_21133), .Q (new_AGEMA_signal_21134) ) ;
    buf_clk new_AGEMA_reg_buffer_8413 ( .C (clk), .D (new_AGEMA_signal_21136), .Q (new_AGEMA_signal_21137) ) ;
    buf_clk new_AGEMA_reg_buffer_8416 ( .C (clk), .D (new_AGEMA_signal_21139), .Q (new_AGEMA_signal_21140) ) ;
    buf_clk new_AGEMA_reg_buffer_8419 ( .C (clk), .D (new_AGEMA_signal_21142), .Q (new_AGEMA_signal_21143) ) ;
    buf_clk new_AGEMA_reg_buffer_8422 ( .C (clk), .D (new_AGEMA_signal_21145), .Q (new_AGEMA_signal_21146) ) ;
    buf_clk new_AGEMA_reg_buffer_8425 ( .C (clk), .D (new_AGEMA_signal_21148), .Q (new_AGEMA_signal_21149) ) ;
    buf_clk new_AGEMA_reg_buffer_8428 ( .C (clk), .D (new_AGEMA_signal_21151), .Q (new_AGEMA_signal_21152) ) ;
    buf_clk new_AGEMA_reg_buffer_8431 ( .C (clk), .D (new_AGEMA_signal_21154), .Q (new_AGEMA_signal_21155) ) ;
    buf_clk new_AGEMA_reg_buffer_8434 ( .C (clk), .D (new_AGEMA_signal_21157), .Q (new_AGEMA_signal_21158) ) ;
    buf_clk new_AGEMA_reg_buffer_8437 ( .C (clk), .D (new_AGEMA_signal_21160), .Q (new_AGEMA_signal_21161) ) ;
    buf_clk new_AGEMA_reg_buffer_8440 ( .C (clk), .D (new_AGEMA_signal_21163), .Q (new_AGEMA_signal_21164) ) ;
    buf_clk new_AGEMA_reg_buffer_8443 ( .C (clk), .D (new_AGEMA_signal_21166), .Q (new_AGEMA_signal_21167) ) ;
    buf_clk new_AGEMA_reg_buffer_8446 ( .C (clk), .D (new_AGEMA_signal_21169), .Q (new_AGEMA_signal_21170) ) ;
    buf_clk new_AGEMA_reg_buffer_8449 ( .C (clk), .D (new_AGEMA_signal_21172), .Q (new_AGEMA_signal_21173) ) ;
    buf_clk new_AGEMA_reg_buffer_8452 ( .C (clk), .D (new_AGEMA_signal_21175), .Q (new_AGEMA_signal_21176) ) ;
    buf_clk new_AGEMA_reg_buffer_8455 ( .C (clk), .D (new_AGEMA_signal_21178), .Q (new_AGEMA_signal_21179) ) ;
    buf_clk new_AGEMA_reg_buffer_8458 ( .C (clk), .D (new_AGEMA_signal_21181), .Q (new_AGEMA_signal_21182) ) ;
    buf_clk new_AGEMA_reg_buffer_8461 ( .C (clk), .D (new_AGEMA_signal_21184), .Q (new_AGEMA_signal_21185) ) ;
    buf_clk new_AGEMA_reg_buffer_8464 ( .C (clk), .D (new_AGEMA_signal_21187), .Q (new_AGEMA_signal_21188) ) ;
    buf_clk new_AGEMA_reg_buffer_8467 ( .C (clk), .D (new_AGEMA_signal_21190), .Q (new_AGEMA_signal_21191) ) ;
    buf_clk new_AGEMA_reg_buffer_8470 ( .C (clk), .D (new_AGEMA_signal_21193), .Q (new_AGEMA_signal_21194) ) ;
    buf_clk new_AGEMA_reg_buffer_8473 ( .C (clk), .D (new_AGEMA_signal_21196), .Q (new_AGEMA_signal_21197) ) ;
    buf_clk new_AGEMA_reg_buffer_8476 ( .C (clk), .D (new_AGEMA_signal_21199), .Q (new_AGEMA_signal_21200) ) ;
    buf_clk new_AGEMA_reg_buffer_8479 ( .C (clk), .D (new_AGEMA_signal_21202), .Q (new_AGEMA_signal_21203) ) ;
    buf_clk new_AGEMA_reg_buffer_8482 ( .C (clk), .D (new_AGEMA_signal_21205), .Q (new_AGEMA_signal_21206) ) ;
    buf_clk new_AGEMA_reg_buffer_8485 ( .C (clk), .D (new_AGEMA_signal_21208), .Q (new_AGEMA_signal_21209) ) ;
    buf_clk new_AGEMA_reg_buffer_8488 ( .C (clk), .D (new_AGEMA_signal_21211), .Q (new_AGEMA_signal_21212) ) ;
    buf_clk new_AGEMA_reg_buffer_8491 ( .C (clk), .D (new_AGEMA_signal_21214), .Q (new_AGEMA_signal_21215) ) ;
    buf_clk new_AGEMA_reg_buffer_8494 ( .C (clk), .D (new_AGEMA_signal_21217), .Q (new_AGEMA_signal_21218) ) ;
    buf_clk new_AGEMA_reg_buffer_8497 ( .C (clk), .D (new_AGEMA_signal_21220), .Q (new_AGEMA_signal_21221) ) ;
    buf_clk new_AGEMA_reg_buffer_8500 ( .C (clk), .D (new_AGEMA_signal_21223), .Q (new_AGEMA_signal_21224) ) ;
    buf_clk new_AGEMA_reg_buffer_8503 ( .C (clk), .D (new_AGEMA_signal_21226), .Q (new_AGEMA_signal_21227) ) ;
    buf_clk new_AGEMA_reg_buffer_8506 ( .C (clk), .D (new_AGEMA_signal_21229), .Q (new_AGEMA_signal_21230) ) ;
    buf_clk new_AGEMA_reg_buffer_8509 ( .C (clk), .D (new_AGEMA_signal_21232), .Q (new_AGEMA_signal_21233) ) ;
    buf_clk new_AGEMA_reg_buffer_8512 ( .C (clk), .D (new_AGEMA_signal_21235), .Q (new_AGEMA_signal_21236) ) ;
    buf_clk new_AGEMA_reg_buffer_8515 ( .C (clk), .D (new_AGEMA_signal_21238), .Q (new_AGEMA_signal_21239) ) ;
    buf_clk new_AGEMA_reg_buffer_8518 ( .C (clk), .D (new_AGEMA_signal_21241), .Q (new_AGEMA_signal_21242) ) ;
    buf_clk new_AGEMA_reg_buffer_8521 ( .C (clk), .D (new_AGEMA_signal_21244), .Q (new_AGEMA_signal_21245) ) ;
    buf_clk new_AGEMA_reg_buffer_8524 ( .C (clk), .D (new_AGEMA_signal_21247), .Q (new_AGEMA_signal_21248) ) ;
    buf_clk new_AGEMA_reg_buffer_8527 ( .C (clk), .D (new_AGEMA_signal_21250), .Q (new_AGEMA_signal_21251) ) ;
    buf_clk new_AGEMA_reg_buffer_8530 ( .C (clk), .D (new_AGEMA_signal_21253), .Q (new_AGEMA_signal_21254) ) ;
    buf_clk new_AGEMA_reg_buffer_8533 ( .C (clk), .D (new_AGEMA_signal_21256), .Q (new_AGEMA_signal_21257) ) ;
    buf_clk new_AGEMA_reg_buffer_8536 ( .C (clk), .D (new_AGEMA_signal_21259), .Q (new_AGEMA_signal_21260) ) ;
    buf_clk new_AGEMA_reg_buffer_8539 ( .C (clk), .D (new_AGEMA_signal_21262), .Q (new_AGEMA_signal_21263) ) ;
    buf_clk new_AGEMA_reg_buffer_8542 ( .C (clk), .D (new_AGEMA_signal_21265), .Q (new_AGEMA_signal_21266) ) ;
    buf_clk new_AGEMA_reg_buffer_8545 ( .C (clk), .D (new_AGEMA_signal_21268), .Q (new_AGEMA_signal_21269) ) ;
    buf_clk new_AGEMA_reg_buffer_8548 ( .C (clk), .D (new_AGEMA_signal_21271), .Q (new_AGEMA_signal_21272) ) ;
    buf_clk new_AGEMA_reg_buffer_8551 ( .C (clk), .D (new_AGEMA_signal_21274), .Q (new_AGEMA_signal_21275) ) ;
    buf_clk new_AGEMA_reg_buffer_8554 ( .C (clk), .D (new_AGEMA_signal_21277), .Q (new_AGEMA_signal_21278) ) ;
    buf_clk new_AGEMA_reg_buffer_8557 ( .C (clk), .D (new_AGEMA_signal_21280), .Q (new_AGEMA_signal_21281) ) ;
    buf_clk new_AGEMA_reg_buffer_8560 ( .C (clk), .D (new_AGEMA_signal_21283), .Q (new_AGEMA_signal_21284) ) ;
    buf_clk new_AGEMA_reg_buffer_8563 ( .C (clk), .D (new_AGEMA_signal_21286), .Q (new_AGEMA_signal_21287) ) ;
    buf_clk new_AGEMA_reg_buffer_8566 ( .C (clk), .D (new_AGEMA_signal_21289), .Q (new_AGEMA_signal_21290) ) ;
    buf_clk new_AGEMA_reg_buffer_8569 ( .C (clk), .D (new_AGEMA_signal_21292), .Q (new_AGEMA_signal_21293) ) ;
    buf_clk new_AGEMA_reg_buffer_8572 ( .C (clk), .D (new_AGEMA_signal_21295), .Q (new_AGEMA_signal_21296) ) ;
    buf_clk new_AGEMA_reg_buffer_8575 ( .C (clk), .D (new_AGEMA_signal_21298), .Q (new_AGEMA_signal_21299) ) ;
    buf_clk new_AGEMA_reg_buffer_8578 ( .C (clk), .D (new_AGEMA_signal_21301), .Q (new_AGEMA_signal_21302) ) ;
    buf_clk new_AGEMA_reg_buffer_8581 ( .C (clk), .D (new_AGEMA_signal_21304), .Q (new_AGEMA_signal_21305) ) ;
    buf_clk new_AGEMA_reg_buffer_8584 ( .C (clk), .D (new_AGEMA_signal_21307), .Q (new_AGEMA_signal_21308) ) ;
    buf_clk new_AGEMA_reg_buffer_8587 ( .C (clk), .D (new_AGEMA_signal_21310), .Q (new_AGEMA_signal_21311) ) ;
    buf_clk new_AGEMA_reg_buffer_8590 ( .C (clk), .D (new_AGEMA_signal_21313), .Q (new_AGEMA_signal_21314) ) ;
    buf_clk new_AGEMA_reg_buffer_8593 ( .C (clk), .D (new_AGEMA_signal_21316), .Q (new_AGEMA_signal_21317) ) ;
    buf_clk new_AGEMA_reg_buffer_8596 ( .C (clk), .D (new_AGEMA_signal_21319), .Q (new_AGEMA_signal_21320) ) ;
    buf_clk new_AGEMA_reg_buffer_8599 ( .C (clk), .D (new_AGEMA_signal_21322), .Q (new_AGEMA_signal_21323) ) ;
    buf_clk new_AGEMA_reg_buffer_8602 ( .C (clk), .D (new_AGEMA_signal_21325), .Q (new_AGEMA_signal_21326) ) ;
    buf_clk new_AGEMA_reg_buffer_8605 ( .C (clk), .D (new_AGEMA_signal_21328), .Q (new_AGEMA_signal_21329) ) ;
    buf_clk new_AGEMA_reg_buffer_8608 ( .C (clk), .D (new_AGEMA_signal_21331), .Q (new_AGEMA_signal_21332) ) ;
    buf_clk new_AGEMA_reg_buffer_8611 ( .C (clk), .D (new_AGEMA_signal_21334), .Q (new_AGEMA_signal_21335) ) ;
    buf_clk new_AGEMA_reg_buffer_8614 ( .C (clk), .D (new_AGEMA_signal_21337), .Q (new_AGEMA_signal_21338) ) ;
    buf_clk new_AGEMA_reg_buffer_8617 ( .C (clk), .D (new_AGEMA_signal_21340), .Q (new_AGEMA_signal_21341) ) ;
    buf_clk new_AGEMA_reg_buffer_8620 ( .C (clk), .D (new_AGEMA_signal_21343), .Q (new_AGEMA_signal_21344) ) ;
    buf_clk new_AGEMA_reg_buffer_8623 ( .C (clk), .D (new_AGEMA_signal_21346), .Q (new_AGEMA_signal_21347) ) ;
    buf_clk new_AGEMA_reg_buffer_8626 ( .C (clk), .D (new_AGEMA_signal_21349), .Q (new_AGEMA_signal_21350) ) ;
    buf_clk new_AGEMA_reg_buffer_8629 ( .C (clk), .D (new_AGEMA_signal_21352), .Q (new_AGEMA_signal_21353) ) ;
    buf_clk new_AGEMA_reg_buffer_8632 ( .C (clk), .D (new_AGEMA_signal_21355), .Q (new_AGEMA_signal_21356) ) ;
    buf_clk new_AGEMA_reg_buffer_8635 ( .C (clk), .D (new_AGEMA_signal_21358), .Q (new_AGEMA_signal_21359) ) ;
    buf_clk new_AGEMA_reg_buffer_8638 ( .C (clk), .D (new_AGEMA_signal_21361), .Q (new_AGEMA_signal_21362) ) ;
    buf_clk new_AGEMA_reg_buffer_8641 ( .C (clk), .D (new_AGEMA_signal_21364), .Q (new_AGEMA_signal_21365) ) ;
    buf_clk new_AGEMA_reg_buffer_8644 ( .C (clk), .D (new_AGEMA_signal_21367), .Q (new_AGEMA_signal_21368) ) ;
    buf_clk new_AGEMA_reg_buffer_8647 ( .C (clk), .D (new_AGEMA_signal_21370), .Q (new_AGEMA_signal_21371) ) ;
    buf_clk new_AGEMA_reg_buffer_8650 ( .C (clk), .D (new_AGEMA_signal_21373), .Q (new_AGEMA_signal_21374) ) ;
    buf_clk new_AGEMA_reg_buffer_8653 ( .C (clk), .D (new_AGEMA_signal_21376), .Q (new_AGEMA_signal_21377) ) ;
    buf_clk new_AGEMA_reg_buffer_8656 ( .C (clk), .D (new_AGEMA_signal_21379), .Q (new_AGEMA_signal_21380) ) ;
    buf_clk new_AGEMA_reg_buffer_8659 ( .C (clk), .D (new_AGEMA_signal_21382), .Q (new_AGEMA_signal_21383) ) ;
    buf_clk new_AGEMA_reg_buffer_8662 ( .C (clk), .D (new_AGEMA_signal_21385), .Q (new_AGEMA_signal_21386) ) ;
    buf_clk new_AGEMA_reg_buffer_8665 ( .C (clk), .D (new_AGEMA_signal_21388), .Q (new_AGEMA_signal_21389) ) ;
    buf_clk new_AGEMA_reg_buffer_8668 ( .C (clk), .D (new_AGEMA_signal_21391), .Q (new_AGEMA_signal_21392) ) ;
    buf_clk new_AGEMA_reg_buffer_8671 ( .C (clk), .D (new_AGEMA_signal_21394), .Q (new_AGEMA_signal_21395) ) ;
    buf_clk new_AGEMA_reg_buffer_8674 ( .C (clk), .D (new_AGEMA_signal_21397), .Q (new_AGEMA_signal_21398) ) ;
    buf_clk new_AGEMA_reg_buffer_8677 ( .C (clk), .D (new_AGEMA_signal_21400), .Q (new_AGEMA_signal_21401) ) ;
    buf_clk new_AGEMA_reg_buffer_8680 ( .C (clk), .D (new_AGEMA_signal_21403), .Q (new_AGEMA_signal_21404) ) ;
    buf_clk new_AGEMA_reg_buffer_8683 ( .C (clk), .D (new_AGEMA_signal_21406), .Q (new_AGEMA_signal_21407) ) ;
    buf_clk new_AGEMA_reg_buffer_8686 ( .C (clk), .D (new_AGEMA_signal_21409), .Q (new_AGEMA_signal_21410) ) ;
    buf_clk new_AGEMA_reg_buffer_8689 ( .C (clk), .D (new_AGEMA_signal_21412), .Q (new_AGEMA_signal_21413) ) ;
    buf_clk new_AGEMA_reg_buffer_8692 ( .C (clk), .D (new_AGEMA_signal_21415), .Q (new_AGEMA_signal_21416) ) ;
    buf_clk new_AGEMA_reg_buffer_8695 ( .C (clk), .D (new_AGEMA_signal_21418), .Q (new_AGEMA_signal_21419) ) ;
    buf_clk new_AGEMA_reg_buffer_8698 ( .C (clk), .D (new_AGEMA_signal_21421), .Q (new_AGEMA_signal_21422) ) ;
    buf_clk new_AGEMA_reg_buffer_8701 ( .C (clk), .D (new_AGEMA_signal_21424), .Q (new_AGEMA_signal_21425) ) ;
    buf_clk new_AGEMA_reg_buffer_8704 ( .C (clk), .D (new_AGEMA_signal_21427), .Q (new_AGEMA_signal_21428) ) ;
    buf_clk new_AGEMA_reg_buffer_8707 ( .C (clk), .D (new_AGEMA_signal_21430), .Q (new_AGEMA_signal_21431) ) ;
    buf_clk new_AGEMA_reg_buffer_8710 ( .C (clk), .D (new_AGEMA_signal_21433), .Q (new_AGEMA_signal_21434) ) ;
    buf_clk new_AGEMA_reg_buffer_8713 ( .C (clk), .D (new_AGEMA_signal_21436), .Q (new_AGEMA_signal_21437) ) ;
    buf_clk new_AGEMA_reg_buffer_8716 ( .C (clk), .D (new_AGEMA_signal_21439), .Q (new_AGEMA_signal_21440) ) ;
    buf_clk new_AGEMA_reg_buffer_8719 ( .C (clk), .D (new_AGEMA_signal_21442), .Q (new_AGEMA_signal_21443) ) ;
    buf_clk new_AGEMA_reg_buffer_8722 ( .C (clk), .D (new_AGEMA_signal_21445), .Q (new_AGEMA_signal_21446) ) ;
    buf_clk new_AGEMA_reg_buffer_8725 ( .C (clk), .D (new_AGEMA_signal_21448), .Q (new_AGEMA_signal_21449) ) ;
    buf_clk new_AGEMA_reg_buffer_8728 ( .C (clk), .D (new_AGEMA_signal_21451), .Q (new_AGEMA_signal_21452) ) ;
    buf_clk new_AGEMA_reg_buffer_8731 ( .C (clk), .D (new_AGEMA_signal_21454), .Q (new_AGEMA_signal_21455) ) ;
    buf_clk new_AGEMA_reg_buffer_8734 ( .C (clk), .D (new_AGEMA_signal_21457), .Q (new_AGEMA_signal_21458) ) ;
    buf_clk new_AGEMA_reg_buffer_8737 ( .C (clk), .D (new_AGEMA_signal_21460), .Q (new_AGEMA_signal_21461) ) ;
    buf_clk new_AGEMA_reg_buffer_8740 ( .C (clk), .D (new_AGEMA_signal_21463), .Q (new_AGEMA_signal_21464) ) ;
    buf_clk new_AGEMA_reg_buffer_8743 ( .C (clk), .D (new_AGEMA_signal_21466), .Q (new_AGEMA_signal_21467) ) ;
    buf_clk new_AGEMA_reg_buffer_8746 ( .C (clk), .D (new_AGEMA_signal_21469), .Q (new_AGEMA_signal_21470) ) ;
    buf_clk new_AGEMA_reg_buffer_8749 ( .C (clk), .D (new_AGEMA_signal_21472), .Q (new_AGEMA_signal_21473) ) ;
    buf_clk new_AGEMA_reg_buffer_8752 ( .C (clk), .D (new_AGEMA_signal_21475), .Q (new_AGEMA_signal_21476) ) ;
    buf_clk new_AGEMA_reg_buffer_8755 ( .C (clk), .D (new_AGEMA_signal_21478), .Q (new_AGEMA_signal_21479) ) ;
    buf_clk new_AGEMA_reg_buffer_8758 ( .C (clk), .D (new_AGEMA_signal_21481), .Q (new_AGEMA_signal_21482) ) ;
    buf_clk new_AGEMA_reg_buffer_8761 ( .C (clk), .D (new_AGEMA_signal_21484), .Q (new_AGEMA_signal_21485) ) ;
    buf_clk new_AGEMA_reg_buffer_8764 ( .C (clk), .D (new_AGEMA_signal_21487), .Q (new_AGEMA_signal_21488) ) ;
    buf_clk new_AGEMA_reg_buffer_8767 ( .C (clk), .D (new_AGEMA_signal_21490), .Q (new_AGEMA_signal_21491) ) ;
    buf_clk new_AGEMA_reg_buffer_8770 ( .C (clk), .D (new_AGEMA_signal_21493), .Q (new_AGEMA_signal_21494) ) ;
    buf_clk new_AGEMA_reg_buffer_8773 ( .C (clk), .D (new_AGEMA_signal_21496), .Q (new_AGEMA_signal_21497) ) ;
    buf_clk new_AGEMA_reg_buffer_8776 ( .C (clk), .D (new_AGEMA_signal_21499), .Q (new_AGEMA_signal_21500) ) ;
    buf_clk new_AGEMA_reg_buffer_8779 ( .C (clk), .D (new_AGEMA_signal_21502), .Q (new_AGEMA_signal_21503) ) ;
    buf_clk new_AGEMA_reg_buffer_8782 ( .C (clk), .D (new_AGEMA_signal_21505), .Q (new_AGEMA_signal_21506) ) ;
    buf_clk new_AGEMA_reg_buffer_8785 ( .C (clk), .D (new_AGEMA_signal_21508), .Q (new_AGEMA_signal_21509) ) ;
    buf_clk new_AGEMA_reg_buffer_8788 ( .C (clk), .D (new_AGEMA_signal_21511), .Q (new_AGEMA_signal_21512) ) ;
    buf_clk new_AGEMA_reg_buffer_8791 ( .C (clk), .D (new_AGEMA_signal_21514), .Q (new_AGEMA_signal_21515) ) ;
    buf_clk new_AGEMA_reg_buffer_8794 ( .C (clk), .D (new_AGEMA_signal_21517), .Q (new_AGEMA_signal_21518) ) ;
    buf_clk new_AGEMA_reg_buffer_8797 ( .C (clk), .D (new_AGEMA_signal_21520), .Q (new_AGEMA_signal_21521) ) ;
    buf_clk new_AGEMA_reg_buffer_8800 ( .C (clk), .D (new_AGEMA_signal_21523), .Q (new_AGEMA_signal_21524) ) ;
    buf_clk new_AGEMA_reg_buffer_8803 ( .C (clk), .D (new_AGEMA_signal_21526), .Q (new_AGEMA_signal_21527) ) ;
    buf_clk new_AGEMA_reg_buffer_8806 ( .C (clk), .D (new_AGEMA_signal_21529), .Q (new_AGEMA_signal_21530) ) ;
    buf_clk new_AGEMA_reg_buffer_8809 ( .C (clk), .D (new_AGEMA_signal_21532), .Q (new_AGEMA_signal_21533) ) ;
    buf_clk new_AGEMA_reg_buffer_8812 ( .C (clk), .D (new_AGEMA_signal_21535), .Q (new_AGEMA_signal_21536) ) ;
    buf_clk new_AGEMA_reg_buffer_8815 ( .C (clk), .D (new_AGEMA_signal_21538), .Q (new_AGEMA_signal_21539) ) ;
    buf_clk new_AGEMA_reg_buffer_8818 ( .C (clk), .D (new_AGEMA_signal_21541), .Q (new_AGEMA_signal_21542) ) ;
    buf_clk new_AGEMA_reg_buffer_8821 ( .C (clk), .D (new_AGEMA_signal_21544), .Q (new_AGEMA_signal_21545) ) ;
    buf_clk new_AGEMA_reg_buffer_8824 ( .C (clk), .D (new_AGEMA_signal_21547), .Q (new_AGEMA_signal_21548) ) ;
    buf_clk new_AGEMA_reg_buffer_8827 ( .C (clk), .D (new_AGEMA_signal_21550), .Q (new_AGEMA_signal_21551) ) ;
    buf_clk new_AGEMA_reg_buffer_8830 ( .C (clk), .D (new_AGEMA_signal_21553), .Q (new_AGEMA_signal_21554) ) ;
    buf_clk new_AGEMA_reg_buffer_8833 ( .C (clk), .D (new_AGEMA_signal_21556), .Q (new_AGEMA_signal_21557) ) ;
    buf_clk new_AGEMA_reg_buffer_8836 ( .C (clk), .D (new_AGEMA_signal_21559), .Q (new_AGEMA_signal_21560) ) ;
    buf_clk new_AGEMA_reg_buffer_8839 ( .C (clk), .D (new_AGEMA_signal_21562), .Q (new_AGEMA_signal_21563) ) ;
    buf_clk new_AGEMA_reg_buffer_8842 ( .C (clk), .D (new_AGEMA_signal_21565), .Q (new_AGEMA_signal_21566) ) ;
    buf_clk new_AGEMA_reg_buffer_8845 ( .C (clk), .D (new_AGEMA_signal_21568), .Q (new_AGEMA_signal_21569) ) ;
    buf_clk new_AGEMA_reg_buffer_8848 ( .C (clk), .D (new_AGEMA_signal_21571), .Q (new_AGEMA_signal_21572) ) ;
    buf_clk new_AGEMA_reg_buffer_8851 ( .C (clk), .D (new_AGEMA_signal_21574), .Q (new_AGEMA_signal_21575) ) ;
    buf_clk new_AGEMA_reg_buffer_8854 ( .C (clk), .D (new_AGEMA_signal_21577), .Q (new_AGEMA_signal_21578) ) ;
    buf_clk new_AGEMA_reg_buffer_8857 ( .C (clk), .D (new_AGEMA_signal_21580), .Q (new_AGEMA_signal_21581) ) ;
    buf_clk new_AGEMA_reg_buffer_8860 ( .C (clk), .D (new_AGEMA_signal_21583), .Q (new_AGEMA_signal_21584) ) ;
    buf_clk new_AGEMA_reg_buffer_8863 ( .C (clk), .D (new_AGEMA_signal_21586), .Q (new_AGEMA_signal_21587) ) ;
    buf_clk new_AGEMA_reg_buffer_8866 ( .C (clk), .D (new_AGEMA_signal_21589), .Q (new_AGEMA_signal_21590) ) ;
    buf_clk new_AGEMA_reg_buffer_8869 ( .C (clk), .D (new_AGEMA_signal_21592), .Q (new_AGEMA_signal_21593) ) ;
    buf_clk new_AGEMA_reg_buffer_8872 ( .C (clk), .D (new_AGEMA_signal_21595), .Q (new_AGEMA_signal_21596) ) ;
    buf_clk new_AGEMA_reg_buffer_8875 ( .C (clk), .D (new_AGEMA_signal_21598), .Q (new_AGEMA_signal_21599) ) ;
    buf_clk new_AGEMA_reg_buffer_8878 ( .C (clk), .D (new_AGEMA_signal_21601), .Q (new_AGEMA_signal_21602) ) ;
    buf_clk new_AGEMA_reg_buffer_8881 ( .C (clk), .D (new_AGEMA_signal_21604), .Q (new_AGEMA_signal_21605) ) ;
    buf_clk new_AGEMA_reg_buffer_8884 ( .C (clk), .D (new_AGEMA_signal_21607), .Q (new_AGEMA_signal_21608) ) ;
    buf_clk new_AGEMA_reg_buffer_8887 ( .C (clk), .D (new_AGEMA_signal_21610), .Q (new_AGEMA_signal_21611) ) ;
    buf_clk new_AGEMA_reg_buffer_8890 ( .C (clk), .D (new_AGEMA_signal_21613), .Q (new_AGEMA_signal_21614) ) ;
    buf_clk new_AGEMA_reg_buffer_8893 ( .C (clk), .D (new_AGEMA_signal_21616), .Q (new_AGEMA_signal_21617) ) ;
    buf_clk new_AGEMA_reg_buffer_8896 ( .C (clk), .D (new_AGEMA_signal_21619), .Q (new_AGEMA_signal_21620) ) ;
    buf_clk new_AGEMA_reg_buffer_8899 ( .C (clk), .D (new_AGEMA_signal_21622), .Q (new_AGEMA_signal_21623) ) ;
    buf_clk new_AGEMA_reg_buffer_8902 ( .C (clk), .D (new_AGEMA_signal_21625), .Q (new_AGEMA_signal_21626) ) ;
    buf_clk new_AGEMA_reg_buffer_8905 ( .C (clk), .D (new_AGEMA_signal_21628), .Q (new_AGEMA_signal_21629) ) ;
    buf_clk new_AGEMA_reg_buffer_8908 ( .C (clk), .D (new_AGEMA_signal_21631), .Q (new_AGEMA_signal_21632) ) ;
    buf_clk new_AGEMA_reg_buffer_8911 ( .C (clk), .D (new_AGEMA_signal_21634), .Q (new_AGEMA_signal_21635) ) ;
    buf_clk new_AGEMA_reg_buffer_8914 ( .C (clk), .D (new_AGEMA_signal_21637), .Q (new_AGEMA_signal_21638) ) ;
    buf_clk new_AGEMA_reg_buffer_8917 ( .C (clk), .D (new_AGEMA_signal_21640), .Q (new_AGEMA_signal_21641) ) ;
    buf_clk new_AGEMA_reg_buffer_8920 ( .C (clk), .D (new_AGEMA_signal_21643), .Q (new_AGEMA_signal_21644) ) ;
    buf_clk new_AGEMA_reg_buffer_8923 ( .C (clk), .D (new_AGEMA_signal_21646), .Q (new_AGEMA_signal_21647) ) ;
    buf_clk new_AGEMA_reg_buffer_8926 ( .C (clk), .D (new_AGEMA_signal_21649), .Q (new_AGEMA_signal_21650) ) ;
    buf_clk new_AGEMA_reg_buffer_8929 ( .C (clk), .D (new_AGEMA_signal_21652), .Q (new_AGEMA_signal_21653) ) ;
    buf_clk new_AGEMA_reg_buffer_8932 ( .C (clk), .D (new_AGEMA_signal_21655), .Q (new_AGEMA_signal_21656) ) ;
    buf_clk new_AGEMA_reg_buffer_8935 ( .C (clk), .D (new_AGEMA_signal_21658), .Q (new_AGEMA_signal_21659) ) ;
    buf_clk new_AGEMA_reg_buffer_8938 ( .C (clk), .D (new_AGEMA_signal_21661), .Q (new_AGEMA_signal_21662) ) ;
    buf_clk new_AGEMA_reg_buffer_8941 ( .C (clk), .D (new_AGEMA_signal_21664), .Q (new_AGEMA_signal_21665) ) ;
    buf_clk new_AGEMA_reg_buffer_8944 ( .C (clk), .D (new_AGEMA_signal_21667), .Q (new_AGEMA_signal_21668) ) ;
    buf_clk new_AGEMA_reg_buffer_8947 ( .C (clk), .D (new_AGEMA_signal_21670), .Q (new_AGEMA_signal_21671) ) ;
    buf_clk new_AGEMA_reg_buffer_8950 ( .C (clk), .D (new_AGEMA_signal_21673), .Q (new_AGEMA_signal_21674) ) ;
    buf_clk new_AGEMA_reg_buffer_8953 ( .C (clk), .D (new_AGEMA_signal_21676), .Q (new_AGEMA_signal_21677) ) ;
    buf_clk new_AGEMA_reg_buffer_8956 ( .C (clk), .D (new_AGEMA_signal_21679), .Q (new_AGEMA_signal_21680) ) ;
    buf_clk new_AGEMA_reg_buffer_8959 ( .C (clk), .D (new_AGEMA_signal_21682), .Q (new_AGEMA_signal_21683) ) ;
    buf_clk new_AGEMA_reg_buffer_8962 ( .C (clk), .D (new_AGEMA_signal_21685), .Q (new_AGEMA_signal_21686) ) ;
    buf_clk new_AGEMA_reg_buffer_8965 ( .C (clk), .D (new_AGEMA_signal_21688), .Q (new_AGEMA_signal_21689) ) ;
    buf_clk new_AGEMA_reg_buffer_8968 ( .C (clk), .D (new_AGEMA_signal_21691), .Q (new_AGEMA_signal_21692) ) ;
    buf_clk new_AGEMA_reg_buffer_8971 ( .C (clk), .D (new_AGEMA_signal_21694), .Q (new_AGEMA_signal_21695) ) ;
    buf_clk new_AGEMA_reg_buffer_8974 ( .C (clk), .D (new_AGEMA_signal_21697), .Q (new_AGEMA_signal_21698) ) ;
    buf_clk new_AGEMA_reg_buffer_8977 ( .C (clk), .D (new_AGEMA_signal_21700), .Q (new_AGEMA_signal_21701) ) ;
    buf_clk new_AGEMA_reg_buffer_8980 ( .C (clk), .D (new_AGEMA_signal_21703), .Q (new_AGEMA_signal_21704) ) ;
    buf_clk new_AGEMA_reg_buffer_8983 ( .C (clk), .D (new_AGEMA_signal_21706), .Q (new_AGEMA_signal_21707) ) ;
    buf_clk new_AGEMA_reg_buffer_8986 ( .C (clk), .D (new_AGEMA_signal_21709), .Q (new_AGEMA_signal_21710) ) ;
    buf_clk new_AGEMA_reg_buffer_8989 ( .C (clk), .D (new_AGEMA_signal_21712), .Q (new_AGEMA_signal_21713) ) ;
    buf_clk new_AGEMA_reg_buffer_8992 ( .C (clk), .D (new_AGEMA_signal_21715), .Q (new_AGEMA_signal_21716) ) ;
    buf_clk new_AGEMA_reg_buffer_8995 ( .C (clk), .D (new_AGEMA_signal_21718), .Q (new_AGEMA_signal_21719) ) ;
    buf_clk new_AGEMA_reg_buffer_8998 ( .C (clk), .D (new_AGEMA_signal_21721), .Q (new_AGEMA_signal_21722) ) ;
    buf_clk new_AGEMA_reg_buffer_9001 ( .C (clk), .D (new_AGEMA_signal_21724), .Q (new_AGEMA_signal_21725) ) ;
    buf_clk new_AGEMA_reg_buffer_9004 ( .C (clk), .D (new_AGEMA_signal_21727), .Q (new_AGEMA_signal_21728) ) ;
    buf_clk new_AGEMA_reg_buffer_9007 ( .C (clk), .D (new_AGEMA_signal_21730), .Q (new_AGEMA_signal_21731) ) ;
    buf_clk new_AGEMA_reg_buffer_9010 ( .C (clk), .D (new_AGEMA_signal_21733), .Q (new_AGEMA_signal_21734) ) ;
    buf_clk new_AGEMA_reg_buffer_9013 ( .C (clk), .D (new_AGEMA_signal_21736), .Q (new_AGEMA_signal_21737) ) ;
    buf_clk new_AGEMA_reg_buffer_9016 ( .C (clk), .D (new_AGEMA_signal_21739), .Q (new_AGEMA_signal_21740) ) ;
    buf_clk new_AGEMA_reg_buffer_9019 ( .C (clk), .D (new_AGEMA_signal_21742), .Q (new_AGEMA_signal_21743) ) ;
    buf_clk new_AGEMA_reg_buffer_9022 ( .C (clk), .D (new_AGEMA_signal_21745), .Q (new_AGEMA_signal_21746) ) ;
    buf_clk new_AGEMA_reg_buffer_9025 ( .C (clk), .D (new_AGEMA_signal_21748), .Q (new_AGEMA_signal_21749) ) ;
    buf_clk new_AGEMA_reg_buffer_9028 ( .C (clk), .D (new_AGEMA_signal_21751), .Q (new_AGEMA_signal_21752) ) ;
    buf_clk new_AGEMA_reg_buffer_9031 ( .C (clk), .D (new_AGEMA_signal_21754), .Q (new_AGEMA_signal_21755) ) ;
    buf_clk new_AGEMA_reg_buffer_9034 ( .C (clk), .D (new_AGEMA_signal_21757), .Q (new_AGEMA_signal_21758) ) ;
    buf_clk new_AGEMA_reg_buffer_9037 ( .C (clk), .D (new_AGEMA_signal_21760), .Q (new_AGEMA_signal_21761) ) ;
    buf_clk new_AGEMA_reg_buffer_9040 ( .C (clk), .D (new_AGEMA_signal_21763), .Q (new_AGEMA_signal_21764) ) ;
    buf_clk new_AGEMA_reg_buffer_9043 ( .C (clk), .D (new_AGEMA_signal_21766), .Q (new_AGEMA_signal_21767) ) ;
    buf_clk new_AGEMA_reg_buffer_9046 ( .C (clk), .D (new_AGEMA_signal_21769), .Q (new_AGEMA_signal_21770) ) ;
    buf_clk new_AGEMA_reg_buffer_9049 ( .C (clk), .D (new_AGEMA_signal_21772), .Q (new_AGEMA_signal_21773) ) ;
    buf_clk new_AGEMA_reg_buffer_9052 ( .C (clk), .D (new_AGEMA_signal_21775), .Q (new_AGEMA_signal_21776) ) ;
    buf_clk new_AGEMA_reg_buffer_9055 ( .C (clk), .D (new_AGEMA_signal_21778), .Q (new_AGEMA_signal_21779) ) ;
    buf_clk new_AGEMA_reg_buffer_9058 ( .C (clk), .D (new_AGEMA_signal_21781), .Q (new_AGEMA_signal_21782) ) ;
    buf_clk new_AGEMA_reg_buffer_9061 ( .C (clk), .D (new_AGEMA_signal_21784), .Q (new_AGEMA_signal_21785) ) ;
    buf_clk new_AGEMA_reg_buffer_9064 ( .C (clk), .D (new_AGEMA_signal_21787), .Q (new_AGEMA_signal_21788) ) ;
    buf_clk new_AGEMA_reg_buffer_9067 ( .C (clk), .D (new_AGEMA_signal_21790), .Q (new_AGEMA_signal_21791) ) ;
    buf_clk new_AGEMA_reg_buffer_9070 ( .C (clk), .D (new_AGEMA_signal_21793), .Q (new_AGEMA_signal_21794) ) ;
    buf_clk new_AGEMA_reg_buffer_9073 ( .C (clk), .D (new_AGEMA_signal_21796), .Q (new_AGEMA_signal_21797) ) ;
    buf_clk new_AGEMA_reg_buffer_9076 ( .C (clk), .D (new_AGEMA_signal_21799), .Q (new_AGEMA_signal_21800) ) ;
    buf_clk new_AGEMA_reg_buffer_9079 ( .C (clk), .D (new_AGEMA_signal_21802), .Q (new_AGEMA_signal_21803) ) ;
    buf_clk new_AGEMA_reg_buffer_9082 ( .C (clk), .D (new_AGEMA_signal_21805), .Q (new_AGEMA_signal_21806) ) ;
    buf_clk new_AGEMA_reg_buffer_9085 ( .C (clk), .D (new_AGEMA_signal_21808), .Q (new_AGEMA_signal_21809) ) ;
    buf_clk new_AGEMA_reg_buffer_9088 ( .C (clk), .D (new_AGEMA_signal_21811), .Q (new_AGEMA_signal_21812) ) ;
    buf_clk new_AGEMA_reg_buffer_9091 ( .C (clk), .D (new_AGEMA_signal_21814), .Q (new_AGEMA_signal_21815) ) ;
    buf_clk new_AGEMA_reg_buffer_9095 ( .C (clk), .D (new_AGEMA_signal_21818), .Q (new_AGEMA_signal_21819) ) ;
    buf_clk new_AGEMA_reg_buffer_9099 ( .C (clk), .D (new_AGEMA_signal_21822), .Q (new_AGEMA_signal_21823) ) ;
    buf_clk new_AGEMA_reg_buffer_9103 ( .C (clk), .D (new_AGEMA_signal_21826), .Q (new_AGEMA_signal_21827) ) ;
    buf_clk new_AGEMA_reg_buffer_9107 ( .C (clk), .D (new_AGEMA_signal_21830), .Q (new_AGEMA_signal_21831) ) ;
    buf_clk new_AGEMA_reg_buffer_9111 ( .C (clk), .D (new_AGEMA_signal_21834), .Q (new_AGEMA_signal_21835) ) ;
    buf_clk new_AGEMA_reg_buffer_9115 ( .C (clk), .D (new_AGEMA_signal_21838), .Q (new_AGEMA_signal_21839) ) ;
    buf_clk new_AGEMA_reg_buffer_9119 ( .C (clk), .D (new_AGEMA_signal_21842), .Q (new_AGEMA_signal_21843) ) ;
    buf_clk new_AGEMA_reg_buffer_9123 ( .C (clk), .D (new_AGEMA_signal_21846), .Q (new_AGEMA_signal_21847) ) ;
    buf_clk new_AGEMA_reg_buffer_9127 ( .C (clk), .D (new_AGEMA_signal_21850), .Q (new_AGEMA_signal_21851) ) ;
    buf_clk new_AGEMA_reg_buffer_9131 ( .C (clk), .D (new_AGEMA_signal_21854), .Q (new_AGEMA_signal_21855) ) ;
    buf_clk new_AGEMA_reg_buffer_9135 ( .C (clk), .D (new_AGEMA_signal_21858), .Q (new_AGEMA_signal_21859) ) ;
    buf_clk new_AGEMA_reg_buffer_9139 ( .C (clk), .D (new_AGEMA_signal_21862), .Q (new_AGEMA_signal_21863) ) ;
    buf_clk new_AGEMA_reg_buffer_9143 ( .C (clk), .D (new_AGEMA_signal_21866), .Q (new_AGEMA_signal_21867) ) ;
    buf_clk new_AGEMA_reg_buffer_9147 ( .C (clk), .D (new_AGEMA_signal_21870), .Q (new_AGEMA_signal_21871) ) ;
    buf_clk new_AGEMA_reg_buffer_9151 ( .C (clk), .D (new_AGEMA_signal_21874), .Q (new_AGEMA_signal_21875) ) ;
    buf_clk new_AGEMA_reg_buffer_9155 ( .C (clk), .D (new_AGEMA_signal_21878), .Q (new_AGEMA_signal_21879) ) ;
    buf_clk new_AGEMA_reg_buffer_9159 ( .C (clk), .D (new_AGEMA_signal_21882), .Q (new_AGEMA_signal_21883) ) ;
    buf_clk new_AGEMA_reg_buffer_9163 ( .C (clk), .D (new_AGEMA_signal_21886), .Q (new_AGEMA_signal_21887) ) ;
    buf_clk new_AGEMA_reg_buffer_9167 ( .C (clk), .D (new_AGEMA_signal_21890), .Q (new_AGEMA_signal_21891) ) ;
    buf_clk new_AGEMA_reg_buffer_9171 ( .C (clk), .D (new_AGEMA_signal_21894), .Q (new_AGEMA_signal_21895) ) ;
    buf_clk new_AGEMA_reg_buffer_9175 ( .C (clk), .D (new_AGEMA_signal_21898), .Q (new_AGEMA_signal_21899) ) ;
    buf_clk new_AGEMA_reg_buffer_9179 ( .C (clk), .D (new_AGEMA_signal_21902), .Q (new_AGEMA_signal_21903) ) ;
    buf_clk new_AGEMA_reg_buffer_9183 ( .C (clk), .D (new_AGEMA_signal_21906), .Q (new_AGEMA_signal_21907) ) ;
    buf_clk new_AGEMA_reg_buffer_9187 ( .C (clk), .D (new_AGEMA_signal_21910), .Q (new_AGEMA_signal_21911) ) ;
    buf_clk new_AGEMA_reg_buffer_9191 ( .C (clk), .D (new_AGEMA_signal_21914), .Q (new_AGEMA_signal_21915) ) ;
    buf_clk new_AGEMA_reg_buffer_9195 ( .C (clk), .D (new_AGEMA_signal_21918), .Q (new_AGEMA_signal_21919) ) ;
    buf_clk new_AGEMA_reg_buffer_9199 ( .C (clk), .D (new_AGEMA_signal_21922), .Q (new_AGEMA_signal_21923) ) ;
    buf_clk new_AGEMA_reg_buffer_9203 ( .C (clk), .D (new_AGEMA_signal_21926), .Q (new_AGEMA_signal_21927) ) ;
    buf_clk new_AGEMA_reg_buffer_9207 ( .C (clk), .D (new_AGEMA_signal_21930), .Q (new_AGEMA_signal_21931) ) ;
    buf_clk new_AGEMA_reg_buffer_9211 ( .C (clk), .D (new_AGEMA_signal_21934), .Q (new_AGEMA_signal_21935) ) ;
    buf_clk new_AGEMA_reg_buffer_9215 ( .C (clk), .D (new_AGEMA_signal_21938), .Q (new_AGEMA_signal_21939) ) ;
    buf_clk new_AGEMA_reg_buffer_9219 ( .C (clk), .D (new_AGEMA_signal_21942), .Q (new_AGEMA_signal_21943) ) ;
    buf_clk new_AGEMA_reg_buffer_9223 ( .C (clk), .D (new_AGEMA_signal_21946), .Q (new_AGEMA_signal_21947) ) ;
    buf_clk new_AGEMA_reg_buffer_9227 ( .C (clk), .D (new_AGEMA_signal_21950), .Q (new_AGEMA_signal_21951) ) ;
    buf_clk new_AGEMA_reg_buffer_9231 ( .C (clk), .D (new_AGEMA_signal_21954), .Q (new_AGEMA_signal_21955) ) ;
    buf_clk new_AGEMA_reg_buffer_9235 ( .C (clk), .D (new_AGEMA_signal_21958), .Q (new_AGEMA_signal_21959) ) ;
    buf_clk new_AGEMA_reg_buffer_9239 ( .C (clk), .D (new_AGEMA_signal_21962), .Q (new_AGEMA_signal_21963) ) ;
    buf_clk new_AGEMA_reg_buffer_9243 ( .C (clk), .D (new_AGEMA_signal_21966), .Q (new_AGEMA_signal_21967) ) ;
    buf_clk new_AGEMA_reg_buffer_9247 ( .C (clk), .D (new_AGEMA_signal_21970), .Q (new_AGEMA_signal_21971) ) ;
    buf_clk new_AGEMA_reg_buffer_9251 ( .C (clk), .D (new_AGEMA_signal_21974), .Q (new_AGEMA_signal_21975) ) ;
    buf_clk new_AGEMA_reg_buffer_9255 ( .C (clk), .D (new_AGEMA_signal_21978), .Q (new_AGEMA_signal_21979) ) ;
    buf_clk new_AGEMA_reg_buffer_9259 ( .C (clk), .D (new_AGEMA_signal_21982), .Q (new_AGEMA_signal_21983) ) ;
    buf_clk new_AGEMA_reg_buffer_9263 ( .C (clk), .D (new_AGEMA_signal_21986), .Q (new_AGEMA_signal_21987) ) ;
    buf_clk new_AGEMA_reg_buffer_9267 ( .C (clk), .D (new_AGEMA_signal_21990), .Q (new_AGEMA_signal_21991) ) ;
    buf_clk new_AGEMA_reg_buffer_9271 ( .C (clk), .D (new_AGEMA_signal_21994), .Q (new_AGEMA_signal_21995) ) ;
    buf_clk new_AGEMA_reg_buffer_9275 ( .C (clk), .D (new_AGEMA_signal_21998), .Q (new_AGEMA_signal_21999) ) ;
    buf_clk new_AGEMA_reg_buffer_9279 ( .C (clk), .D (new_AGEMA_signal_22002), .Q (new_AGEMA_signal_22003) ) ;
    buf_clk new_AGEMA_reg_buffer_9283 ( .C (clk), .D (new_AGEMA_signal_22006), .Q (new_AGEMA_signal_22007) ) ;
    buf_clk new_AGEMA_reg_buffer_9287 ( .C (clk), .D (new_AGEMA_signal_22010), .Q (new_AGEMA_signal_22011) ) ;
    buf_clk new_AGEMA_reg_buffer_9291 ( .C (clk), .D (new_AGEMA_signal_22014), .Q (new_AGEMA_signal_22015) ) ;
    buf_clk new_AGEMA_reg_buffer_9295 ( .C (clk), .D (new_AGEMA_signal_22018), .Q (new_AGEMA_signal_22019) ) ;
    buf_clk new_AGEMA_reg_buffer_9299 ( .C (clk), .D (new_AGEMA_signal_22022), .Q (new_AGEMA_signal_22023) ) ;
    buf_clk new_AGEMA_reg_buffer_9303 ( .C (clk), .D (new_AGEMA_signal_22026), .Q (new_AGEMA_signal_22027) ) ;
    buf_clk new_AGEMA_reg_buffer_9307 ( .C (clk), .D (new_AGEMA_signal_22030), .Q (new_AGEMA_signal_22031) ) ;
    buf_clk new_AGEMA_reg_buffer_9311 ( .C (clk), .D (new_AGEMA_signal_22034), .Q (new_AGEMA_signal_22035) ) ;
    buf_clk new_AGEMA_reg_buffer_9315 ( .C (clk), .D (new_AGEMA_signal_22038), .Q (new_AGEMA_signal_22039) ) ;
    buf_clk new_AGEMA_reg_buffer_9319 ( .C (clk), .D (new_AGEMA_signal_22042), .Q (new_AGEMA_signal_22043) ) ;
    buf_clk new_AGEMA_reg_buffer_9323 ( .C (clk), .D (new_AGEMA_signal_22046), .Q (new_AGEMA_signal_22047) ) ;
    buf_clk new_AGEMA_reg_buffer_9327 ( .C (clk), .D (new_AGEMA_signal_22050), .Q (new_AGEMA_signal_22051) ) ;
    buf_clk new_AGEMA_reg_buffer_9331 ( .C (clk), .D (new_AGEMA_signal_22054), .Q (new_AGEMA_signal_22055) ) ;
    buf_clk new_AGEMA_reg_buffer_9335 ( .C (clk), .D (new_AGEMA_signal_22058), .Q (new_AGEMA_signal_22059) ) ;
    buf_clk new_AGEMA_reg_buffer_9339 ( .C (clk), .D (new_AGEMA_signal_22062), .Q (new_AGEMA_signal_22063) ) ;
    buf_clk new_AGEMA_reg_buffer_9343 ( .C (clk), .D (new_AGEMA_signal_22066), .Q (new_AGEMA_signal_22067) ) ;
    buf_clk new_AGEMA_reg_buffer_9347 ( .C (clk), .D (new_AGEMA_signal_22070), .Q (new_AGEMA_signal_22071) ) ;
    buf_clk new_AGEMA_reg_buffer_9351 ( .C (clk), .D (new_AGEMA_signal_22074), .Q (new_AGEMA_signal_22075) ) ;
    buf_clk new_AGEMA_reg_buffer_9355 ( .C (clk), .D (new_AGEMA_signal_22078), .Q (new_AGEMA_signal_22079) ) ;
    buf_clk new_AGEMA_reg_buffer_9359 ( .C (clk), .D (new_AGEMA_signal_22082), .Q (new_AGEMA_signal_22083) ) ;
    buf_clk new_AGEMA_reg_buffer_9363 ( .C (clk), .D (new_AGEMA_signal_22086), .Q (new_AGEMA_signal_22087) ) ;
    buf_clk new_AGEMA_reg_buffer_9367 ( .C (clk), .D (new_AGEMA_signal_22090), .Q (new_AGEMA_signal_22091) ) ;
    buf_clk new_AGEMA_reg_buffer_9371 ( .C (clk), .D (new_AGEMA_signal_22094), .Q (new_AGEMA_signal_22095) ) ;
    buf_clk new_AGEMA_reg_buffer_9375 ( .C (clk), .D (new_AGEMA_signal_22098), .Q (new_AGEMA_signal_22099) ) ;
    buf_clk new_AGEMA_reg_buffer_9379 ( .C (clk), .D (new_AGEMA_signal_22102), .Q (new_AGEMA_signal_22103) ) ;
    buf_clk new_AGEMA_reg_buffer_9383 ( .C (clk), .D (new_AGEMA_signal_22106), .Q (new_AGEMA_signal_22107) ) ;
    buf_clk new_AGEMA_reg_buffer_9387 ( .C (clk), .D (new_AGEMA_signal_22110), .Q (new_AGEMA_signal_22111) ) ;
    buf_clk new_AGEMA_reg_buffer_9391 ( .C (clk), .D (new_AGEMA_signal_22114), .Q (new_AGEMA_signal_22115) ) ;
    buf_clk new_AGEMA_reg_buffer_9395 ( .C (clk), .D (new_AGEMA_signal_22118), .Q (new_AGEMA_signal_22119) ) ;
    buf_clk new_AGEMA_reg_buffer_9399 ( .C (clk), .D (new_AGEMA_signal_22122), .Q (new_AGEMA_signal_22123) ) ;
    buf_clk new_AGEMA_reg_buffer_9403 ( .C (clk), .D (new_AGEMA_signal_22126), .Q (new_AGEMA_signal_22127) ) ;
    buf_clk new_AGEMA_reg_buffer_9407 ( .C (clk), .D (new_AGEMA_signal_22130), .Q (new_AGEMA_signal_22131) ) ;
    buf_clk new_AGEMA_reg_buffer_9411 ( .C (clk), .D (new_AGEMA_signal_22134), .Q (new_AGEMA_signal_22135) ) ;
    buf_clk new_AGEMA_reg_buffer_9415 ( .C (clk), .D (new_AGEMA_signal_22138), .Q (new_AGEMA_signal_22139) ) ;
    buf_clk new_AGEMA_reg_buffer_9419 ( .C (clk), .D (new_AGEMA_signal_22142), .Q (new_AGEMA_signal_22143) ) ;
    buf_clk new_AGEMA_reg_buffer_9423 ( .C (clk), .D (new_AGEMA_signal_22146), .Q (new_AGEMA_signal_22147) ) ;
    buf_clk new_AGEMA_reg_buffer_9427 ( .C (clk), .D (new_AGEMA_signal_22150), .Q (new_AGEMA_signal_22151) ) ;
    buf_clk new_AGEMA_reg_buffer_9431 ( .C (clk), .D (new_AGEMA_signal_22154), .Q (new_AGEMA_signal_22155) ) ;
    buf_clk new_AGEMA_reg_buffer_9435 ( .C (clk), .D (new_AGEMA_signal_22158), .Q (new_AGEMA_signal_22159) ) ;
    buf_clk new_AGEMA_reg_buffer_9439 ( .C (clk), .D (new_AGEMA_signal_22162), .Q (new_AGEMA_signal_22163) ) ;
    buf_clk new_AGEMA_reg_buffer_9443 ( .C (clk), .D (new_AGEMA_signal_22166), .Q (new_AGEMA_signal_22167) ) ;
    buf_clk new_AGEMA_reg_buffer_9447 ( .C (clk), .D (new_AGEMA_signal_22170), .Q (new_AGEMA_signal_22171) ) ;
    buf_clk new_AGEMA_reg_buffer_9451 ( .C (clk), .D (new_AGEMA_signal_22174), .Q (new_AGEMA_signal_22175) ) ;
    buf_clk new_AGEMA_reg_buffer_9455 ( .C (clk), .D (new_AGEMA_signal_22178), .Q (new_AGEMA_signal_22179) ) ;
    buf_clk new_AGEMA_reg_buffer_9459 ( .C (clk), .D (new_AGEMA_signal_22182), .Q (new_AGEMA_signal_22183) ) ;
    buf_clk new_AGEMA_reg_buffer_9463 ( .C (clk), .D (new_AGEMA_signal_22186), .Q (new_AGEMA_signal_22187) ) ;
    buf_clk new_AGEMA_reg_buffer_9467 ( .C (clk), .D (new_AGEMA_signal_22190), .Q (new_AGEMA_signal_22191) ) ;
    buf_clk new_AGEMA_reg_buffer_9471 ( .C (clk), .D (new_AGEMA_signal_22194), .Q (new_AGEMA_signal_22195) ) ;
    buf_clk new_AGEMA_reg_buffer_9475 ( .C (clk), .D (new_AGEMA_signal_22198), .Q (new_AGEMA_signal_22199) ) ;
    buf_clk new_AGEMA_reg_buffer_9479 ( .C (clk), .D (new_AGEMA_signal_22202), .Q (new_AGEMA_signal_22203) ) ;
    buf_clk new_AGEMA_reg_buffer_9483 ( .C (clk), .D (new_AGEMA_signal_22206), .Q (new_AGEMA_signal_22207) ) ;
    buf_clk new_AGEMA_reg_buffer_9487 ( .C (clk), .D (new_AGEMA_signal_22210), .Q (new_AGEMA_signal_22211) ) ;
    buf_clk new_AGEMA_reg_buffer_9491 ( .C (clk), .D (new_AGEMA_signal_22214), .Q (new_AGEMA_signal_22215) ) ;
    buf_clk new_AGEMA_reg_buffer_9495 ( .C (clk), .D (new_AGEMA_signal_22218), .Q (new_AGEMA_signal_22219) ) ;
    buf_clk new_AGEMA_reg_buffer_9499 ( .C (clk), .D (new_AGEMA_signal_22222), .Q (new_AGEMA_signal_22223) ) ;
    buf_clk new_AGEMA_reg_buffer_9503 ( .C (clk), .D (new_AGEMA_signal_22226), .Q (new_AGEMA_signal_22227) ) ;
    buf_clk new_AGEMA_reg_buffer_9507 ( .C (clk), .D (new_AGEMA_signal_22230), .Q (new_AGEMA_signal_22231) ) ;
    buf_clk new_AGEMA_reg_buffer_9511 ( .C (clk), .D (new_AGEMA_signal_22234), .Q (new_AGEMA_signal_22235) ) ;
    buf_clk new_AGEMA_reg_buffer_9515 ( .C (clk), .D (new_AGEMA_signal_22238), .Q (new_AGEMA_signal_22239) ) ;
    buf_clk new_AGEMA_reg_buffer_9519 ( .C (clk), .D (new_AGEMA_signal_22242), .Q (new_AGEMA_signal_22243) ) ;
    buf_clk new_AGEMA_reg_buffer_9523 ( .C (clk), .D (new_AGEMA_signal_22246), .Q (new_AGEMA_signal_22247) ) ;
    buf_clk new_AGEMA_reg_buffer_9527 ( .C (clk), .D (new_AGEMA_signal_22250), .Q (new_AGEMA_signal_22251) ) ;
    buf_clk new_AGEMA_reg_buffer_9531 ( .C (clk), .D (new_AGEMA_signal_22254), .Q (new_AGEMA_signal_22255) ) ;
    buf_clk new_AGEMA_reg_buffer_9535 ( .C (clk), .D (new_AGEMA_signal_22258), .Q (new_AGEMA_signal_22259) ) ;
    buf_clk new_AGEMA_reg_buffer_9539 ( .C (clk), .D (new_AGEMA_signal_22262), .Q (new_AGEMA_signal_22263) ) ;
    buf_clk new_AGEMA_reg_buffer_9543 ( .C (clk), .D (new_AGEMA_signal_22266), .Q (new_AGEMA_signal_22267) ) ;
    buf_clk new_AGEMA_reg_buffer_9547 ( .C (clk), .D (new_AGEMA_signal_22270), .Q (new_AGEMA_signal_22271) ) ;
    buf_clk new_AGEMA_reg_buffer_9551 ( .C (clk), .D (new_AGEMA_signal_22274), .Q (new_AGEMA_signal_22275) ) ;
    buf_clk new_AGEMA_reg_buffer_9555 ( .C (clk), .D (new_AGEMA_signal_22278), .Q (new_AGEMA_signal_22279) ) ;
    buf_clk new_AGEMA_reg_buffer_9559 ( .C (clk), .D (new_AGEMA_signal_22282), .Q (new_AGEMA_signal_22283) ) ;
    buf_clk new_AGEMA_reg_buffer_9563 ( .C (clk), .D (new_AGEMA_signal_22286), .Q (new_AGEMA_signal_22287) ) ;
    buf_clk new_AGEMA_reg_buffer_9567 ( .C (clk), .D (new_AGEMA_signal_22290), .Q (new_AGEMA_signal_22291) ) ;
    buf_clk new_AGEMA_reg_buffer_9571 ( .C (clk), .D (new_AGEMA_signal_22294), .Q (new_AGEMA_signal_22295) ) ;
    buf_clk new_AGEMA_reg_buffer_9575 ( .C (clk), .D (new_AGEMA_signal_22298), .Q (new_AGEMA_signal_22299) ) ;
    buf_clk new_AGEMA_reg_buffer_9579 ( .C (clk), .D (new_AGEMA_signal_22302), .Q (new_AGEMA_signal_22303) ) ;
    buf_clk new_AGEMA_reg_buffer_9583 ( .C (clk), .D (new_AGEMA_signal_22306), .Q (new_AGEMA_signal_22307) ) ;
    buf_clk new_AGEMA_reg_buffer_9587 ( .C (clk), .D (new_AGEMA_signal_22310), .Q (new_AGEMA_signal_22311) ) ;
    buf_clk new_AGEMA_reg_buffer_9591 ( .C (clk), .D (new_AGEMA_signal_22314), .Q (new_AGEMA_signal_22315) ) ;
    buf_clk new_AGEMA_reg_buffer_9595 ( .C (clk), .D (new_AGEMA_signal_22318), .Q (new_AGEMA_signal_22319) ) ;
    buf_clk new_AGEMA_reg_buffer_9599 ( .C (clk), .D (new_AGEMA_signal_22322), .Q (new_AGEMA_signal_22323) ) ;
    buf_clk new_AGEMA_reg_buffer_9603 ( .C (clk), .D (new_AGEMA_signal_22326), .Q (new_AGEMA_signal_22327) ) ;
    buf_clk new_AGEMA_reg_buffer_9607 ( .C (clk), .D (new_AGEMA_signal_22330), .Q (new_AGEMA_signal_22331) ) ;
    buf_clk new_AGEMA_reg_buffer_9611 ( .C (clk), .D (new_AGEMA_signal_22334), .Q (new_AGEMA_signal_22335) ) ;
    buf_clk new_AGEMA_reg_buffer_9615 ( .C (clk), .D (new_AGEMA_signal_22338), .Q (new_AGEMA_signal_22339) ) ;
    buf_clk new_AGEMA_reg_buffer_9619 ( .C (clk), .D (new_AGEMA_signal_22342), .Q (new_AGEMA_signal_22343) ) ;
    buf_clk new_AGEMA_reg_buffer_9623 ( .C (clk), .D (new_AGEMA_signal_22346), .Q (new_AGEMA_signal_22347) ) ;
    buf_clk new_AGEMA_reg_buffer_9627 ( .C (clk), .D (new_AGEMA_signal_22350), .Q (new_AGEMA_signal_22351) ) ;
    buf_clk new_AGEMA_reg_buffer_9631 ( .C (clk), .D (new_AGEMA_signal_22354), .Q (new_AGEMA_signal_22355) ) ;
    buf_clk new_AGEMA_reg_buffer_9635 ( .C (clk), .D (new_AGEMA_signal_22358), .Q (new_AGEMA_signal_22359) ) ;
    buf_clk new_AGEMA_reg_buffer_9639 ( .C (clk), .D (new_AGEMA_signal_22362), .Q (new_AGEMA_signal_22363) ) ;
    buf_clk new_AGEMA_reg_buffer_9643 ( .C (clk), .D (new_AGEMA_signal_22366), .Q (new_AGEMA_signal_22367) ) ;
    buf_clk new_AGEMA_reg_buffer_9647 ( .C (clk), .D (new_AGEMA_signal_22370), .Q (new_AGEMA_signal_22371) ) ;
    buf_clk new_AGEMA_reg_buffer_9651 ( .C (clk), .D (new_AGEMA_signal_22374), .Q (new_AGEMA_signal_22375) ) ;
    buf_clk new_AGEMA_reg_buffer_9655 ( .C (clk), .D (new_AGEMA_signal_22378), .Q (new_AGEMA_signal_22379) ) ;
    buf_clk new_AGEMA_reg_buffer_9659 ( .C (clk), .D (new_AGEMA_signal_22382), .Q (new_AGEMA_signal_22383) ) ;
    buf_clk new_AGEMA_reg_buffer_9663 ( .C (clk), .D (new_AGEMA_signal_22386), .Q (new_AGEMA_signal_22387) ) ;
    buf_clk new_AGEMA_reg_buffer_9667 ( .C (clk), .D (new_AGEMA_signal_22390), .Q (new_AGEMA_signal_22391) ) ;
    buf_clk new_AGEMA_reg_buffer_9671 ( .C (clk), .D (new_AGEMA_signal_22394), .Q (new_AGEMA_signal_22395) ) ;
    buf_clk new_AGEMA_reg_buffer_9675 ( .C (clk), .D (new_AGEMA_signal_22398), .Q (new_AGEMA_signal_22399) ) ;
    buf_clk new_AGEMA_reg_buffer_9679 ( .C (clk), .D (new_AGEMA_signal_22402), .Q (new_AGEMA_signal_22403) ) ;
    buf_clk new_AGEMA_reg_buffer_9683 ( .C (clk), .D (new_AGEMA_signal_22406), .Q (new_AGEMA_signal_22407) ) ;
    buf_clk new_AGEMA_reg_buffer_9687 ( .C (clk), .D (new_AGEMA_signal_22410), .Q (new_AGEMA_signal_22411) ) ;
    buf_clk new_AGEMA_reg_buffer_9691 ( .C (clk), .D (new_AGEMA_signal_22414), .Q (new_AGEMA_signal_22415) ) ;
    buf_clk new_AGEMA_reg_buffer_9695 ( .C (clk), .D (new_AGEMA_signal_22418), .Q (new_AGEMA_signal_22419) ) ;
    buf_clk new_AGEMA_reg_buffer_9699 ( .C (clk), .D (new_AGEMA_signal_22422), .Q (new_AGEMA_signal_22423) ) ;
    buf_clk new_AGEMA_reg_buffer_9703 ( .C (clk), .D (new_AGEMA_signal_22426), .Q (new_AGEMA_signal_22427) ) ;
    buf_clk new_AGEMA_reg_buffer_9707 ( .C (clk), .D (new_AGEMA_signal_22430), .Q (new_AGEMA_signal_22431) ) ;
    buf_clk new_AGEMA_reg_buffer_9711 ( .C (clk), .D (new_AGEMA_signal_22434), .Q (new_AGEMA_signal_22435) ) ;
    buf_clk new_AGEMA_reg_buffer_9715 ( .C (clk), .D (new_AGEMA_signal_22438), .Q (new_AGEMA_signal_22439) ) ;
    buf_clk new_AGEMA_reg_buffer_9719 ( .C (clk), .D (new_AGEMA_signal_22442), .Q (new_AGEMA_signal_22443) ) ;
    buf_clk new_AGEMA_reg_buffer_9723 ( .C (clk), .D (new_AGEMA_signal_22446), .Q (new_AGEMA_signal_22447) ) ;
    buf_clk new_AGEMA_reg_buffer_9727 ( .C (clk), .D (new_AGEMA_signal_22450), .Q (new_AGEMA_signal_22451) ) ;
    buf_clk new_AGEMA_reg_buffer_9731 ( .C (clk), .D (new_AGEMA_signal_22454), .Q (new_AGEMA_signal_22455) ) ;
    buf_clk new_AGEMA_reg_buffer_9735 ( .C (clk), .D (new_AGEMA_signal_22458), .Q (new_AGEMA_signal_22459) ) ;
    buf_clk new_AGEMA_reg_buffer_9739 ( .C (clk), .D (new_AGEMA_signal_22462), .Q (new_AGEMA_signal_22463) ) ;
    buf_clk new_AGEMA_reg_buffer_9743 ( .C (clk), .D (new_AGEMA_signal_22466), .Q (new_AGEMA_signal_22467) ) ;
    buf_clk new_AGEMA_reg_buffer_9747 ( .C (clk), .D (new_AGEMA_signal_22470), .Q (new_AGEMA_signal_22471) ) ;
    buf_clk new_AGEMA_reg_buffer_9751 ( .C (clk), .D (new_AGEMA_signal_22474), .Q (new_AGEMA_signal_22475) ) ;
    buf_clk new_AGEMA_reg_buffer_9755 ( .C (clk), .D (new_AGEMA_signal_22478), .Q (new_AGEMA_signal_22479) ) ;
    buf_clk new_AGEMA_reg_buffer_9759 ( .C (clk), .D (new_AGEMA_signal_22482), .Q (new_AGEMA_signal_22483) ) ;
    buf_clk new_AGEMA_reg_buffer_9763 ( .C (clk), .D (new_AGEMA_signal_22486), .Q (new_AGEMA_signal_22487) ) ;
    buf_clk new_AGEMA_reg_buffer_9767 ( .C (clk), .D (new_AGEMA_signal_22490), .Q (new_AGEMA_signal_22491) ) ;
    buf_clk new_AGEMA_reg_buffer_9771 ( .C (clk), .D (new_AGEMA_signal_22494), .Q (new_AGEMA_signal_22495) ) ;
    buf_clk new_AGEMA_reg_buffer_9775 ( .C (clk), .D (new_AGEMA_signal_22498), .Q (new_AGEMA_signal_22499) ) ;
    buf_clk new_AGEMA_reg_buffer_9779 ( .C (clk), .D (new_AGEMA_signal_22502), .Q (new_AGEMA_signal_22503) ) ;
    buf_clk new_AGEMA_reg_buffer_9783 ( .C (clk), .D (new_AGEMA_signal_22506), .Q (new_AGEMA_signal_22507) ) ;
    buf_clk new_AGEMA_reg_buffer_9787 ( .C (clk), .D (new_AGEMA_signal_22510), .Q (new_AGEMA_signal_22511) ) ;
    buf_clk new_AGEMA_reg_buffer_9791 ( .C (clk), .D (new_AGEMA_signal_22514), .Q (new_AGEMA_signal_22515) ) ;
    buf_clk new_AGEMA_reg_buffer_9795 ( .C (clk), .D (new_AGEMA_signal_22518), .Q (new_AGEMA_signal_22519) ) ;
    buf_clk new_AGEMA_reg_buffer_9799 ( .C (clk), .D (new_AGEMA_signal_22522), .Q (new_AGEMA_signal_22523) ) ;
    buf_clk new_AGEMA_reg_buffer_9803 ( .C (clk), .D (new_AGEMA_signal_22526), .Q (new_AGEMA_signal_22527) ) ;
    buf_clk new_AGEMA_reg_buffer_9807 ( .C (clk), .D (new_AGEMA_signal_22530), .Q (new_AGEMA_signal_22531) ) ;
    buf_clk new_AGEMA_reg_buffer_9811 ( .C (clk), .D (new_AGEMA_signal_22534), .Q (new_AGEMA_signal_22535) ) ;
    buf_clk new_AGEMA_reg_buffer_9815 ( .C (clk), .D (new_AGEMA_signal_22538), .Q (new_AGEMA_signal_22539) ) ;
    buf_clk new_AGEMA_reg_buffer_9819 ( .C (clk), .D (new_AGEMA_signal_22542), .Q (new_AGEMA_signal_22543) ) ;
    buf_clk new_AGEMA_reg_buffer_9823 ( .C (clk), .D (new_AGEMA_signal_22546), .Q (new_AGEMA_signal_22547) ) ;
    buf_clk new_AGEMA_reg_buffer_9827 ( .C (clk), .D (new_AGEMA_signal_22550), .Q (new_AGEMA_signal_22551) ) ;
    buf_clk new_AGEMA_reg_buffer_9831 ( .C (clk), .D (new_AGEMA_signal_22554), .Q (new_AGEMA_signal_22555) ) ;
    buf_clk new_AGEMA_reg_buffer_9835 ( .C (clk), .D (new_AGEMA_signal_22558), .Q (new_AGEMA_signal_22559) ) ;
    buf_clk new_AGEMA_reg_buffer_9839 ( .C (clk), .D (new_AGEMA_signal_22562), .Q (new_AGEMA_signal_22563) ) ;
    buf_clk new_AGEMA_reg_buffer_9843 ( .C (clk), .D (new_AGEMA_signal_22566), .Q (new_AGEMA_signal_22567) ) ;
    buf_clk new_AGEMA_reg_buffer_9847 ( .C (clk), .D (new_AGEMA_signal_22570), .Q (new_AGEMA_signal_22571) ) ;
    buf_clk new_AGEMA_reg_buffer_9851 ( .C (clk), .D (new_AGEMA_signal_22574), .Q (new_AGEMA_signal_22575) ) ;
    buf_clk new_AGEMA_reg_buffer_9855 ( .C (clk), .D (new_AGEMA_signal_22578), .Q (new_AGEMA_signal_22579) ) ;
    buf_clk new_AGEMA_reg_buffer_9859 ( .C (clk), .D (new_AGEMA_signal_22582), .Q (new_AGEMA_signal_22583) ) ;
    buf_clk new_AGEMA_reg_buffer_9863 ( .C (clk), .D (new_AGEMA_signal_22586), .Q (new_AGEMA_signal_22587) ) ;
    buf_clk new_AGEMA_reg_buffer_9867 ( .C (clk), .D (new_AGEMA_signal_22590), .Q (new_AGEMA_signal_22591) ) ;
    buf_clk new_AGEMA_reg_buffer_9871 ( .C (clk), .D (new_AGEMA_signal_22594), .Q (new_AGEMA_signal_22595) ) ;
    buf_clk new_AGEMA_reg_buffer_9875 ( .C (clk), .D (new_AGEMA_signal_22598), .Q (new_AGEMA_signal_22599) ) ;
    buf_clk new_AGEMA_reg_buffer_9879 ( .C (clk), .D (new_AGEMA_signal_22602), .Q (new_AGEMA_signal_22603) ) ;
    buf_clk new_AGEMA_reg_buffer_9883 ( .C (clk), .D (new_AGEMA_signal_22606), .Q (new_AGEMA_signal_22607) ) ;
    buf_clk new_AGEMA_reg_buffer_9887 ( .C (clk), .D (new_AGEMA_signal_22610), .Q (new_AGEMA_signal_22611) ) ;
    buf_clk new_AGEMA_reg_buffer_9891 ( .C (clk), .D (new_AGEMA_signal_22614), .Q (new_AGEMA_signal_22615) ) ;
    buf_clk new_AGEMA_reg_buffer_9895 ( .C (clk), .D (new_AGEMA_signal_22618), .Q (new_AGEMA_signal_22619) ) ;
    buf_clk new_AGEMA_reg_buffer_9899 ( .C (clk), .D (new_AGEMA_signal_22622), .Q (new_AGEMA_signal_22623) ) ;
    buf_clk new_AGEMA_reg_buffer_9903 ( .C (clk), .D (new_AGEMA_signal_22626), .Q (new_AGEMA_signal_22627) ) ;
    buf_clk new_AGEMA_reg_buffer_9907 ( .C (clk), .D (new_AGEMA_signal_22630), .Q (new_AGEMA_signal_22631) ) ;
    buf_clk new_AGEMA_reg_buffer_9911 ( .C (clk), .D (new_AGEMA_signal_22634), .Q (new_AGEMA_signal_22635) ) ;
    buf_clk new_AGEMA_reg_buffer_9915 ( .C (clk), .D (new_AGEMA_signal_22638), .Q (new_AGEMA_signal_22639) ) ;
    buf_clk new_AGEMA_reg_buffer_9919 ( .C (clk), .D (new_AGEMA_signal_22642), .Q (new_AGEMA_signal_22643) ) ;
    buf_clk new_AGEMA_reg_buffer_9923 ( .C (clk), .D (new_AGEMA_signal_22646), .Q (new_AGEMA_signal_22647) ) ;
    buf_clk new_AGEMA_reg_buffer_9927 ( .C (clk), .D (new_AGEMA_signal_22650), .Q (new_AGEMA_signal_22651) ) ;
    buf_clk new_AGEMA_reg_buffer_9931 ( .C (clk), .D (new_AGEMA_signal_22654), .Q (new_AGEMA_signal_22655) ) ;
    buf_clk new_AGEMA_reg_buffer_9935 ( .C (clk), .D (new_AGEMA_signal_22658), .Q (new_AGEMA_signal_22659) ) ;
    buf_clk new_AGEMA_reg_buffer_9939 ( .C (clk), .D (new_AGEMA_signal_22662), .Q (new_AGEMA_signal_22663) ) ;
    buf_clk new_AGEMA_reg_buffer_9943 ( .C (clk), .D (new_AGEMA_signal_22666), .Q (new_AGEMA_signal_22667) ) ;
    buf_clk new_AGEMA_reg_buffer_9947 ( .C (clk), .D (new_AGEMA_signal_22670), .Q (new_AGEMA_signal_22671) ) ;
    buf_clk new_AGEMA_reg_buffer_9951 ( .C (clk), .D (new_AGEMA_signal_22674), .Q (new_AGEMA_signal_22675) ) ;
    buf_clk new_AGEMA_reg_buffer_9955 ( .C (clk), .D (new_AGEMA_signal_22678), .Q (new_AGEMA_signal_22679) ) ;
    buf_clk new_AGEMA_reg_buffer_9959 ( .C (clk), .D (new_AGEMA_signal_22682), .Q (new_AGEMA_signal_22683) ) ;
    buf_clk new_AGEMA_reg_buffer_9963 ( .C (clk), .D (new_AGEMA_signal_22686), .Q (new_AGEMA_signal_22687) ) ;
    buf_clk new_AGEMA_reg_buffer_9967 ( .C (clk), .D (new_AGEMA_signal_22690), .Q (new_AGEMA_signal_22691) ) ;
    buf_clk new_AGEMA_reg_buffer_9971 ( .C (clk), .D (new_AGEMA_signal_22694), .Q (new_AGEMA_signal_22695) ) ;
    buf_clk new_AGEMA_reg_buffer_9975 ( .C (clk), .D (new_AGEMA_signal_22698), .Q (new_AGEMA_signal_22699) ) ;
    buf_clk new_AGEMA_reg_buffer_9979 ( .C (clk), .D (new_AGEMA_signal_22702), .Q (new_AGEMA_signal_22703) ) ;
    buf_clk new_AGEMA_reg_buffer_9983 ( .C (clk), .D (new_AGEMA_signal_22706), .Q (new_AGEMA_signal_22707) ) ;
    buf_clk new_AGEMA_reg_buffer_9987 ( .C (clk), .D (new_AGEMA_signal_22710), .Q (new_AGEMA_signal_22711) ) ;
    buf_clk new_AGEMA_reg_buffer_9991 ( .C (clk), .D (new_AGEMA_signal_22714), .Q (new_AGEMA_signal_22715) ) ;
    buf_clk new_AGEMA_reg_buffer_9995 ( .C (clk), .D (new_AGEMA_signal_22718), .Q (new_AGEMA_signal_22719) ) ;
    buf_clk new_AGEMA_reg_buffer_9999 ( .C (clk), .D (new_AGEMA_signal_22722), .Q (new_AGEMA_signal_22723) ) ;
    buf_clk new_AGEMA_reg_buffer_10003 ( .C (clk), .D (new_AGEMA_signal_22726), .Q (new_AGEMA_signal_22727) ) ;
    buf_clk new_AGEMA_reg_buffer_10007 ( .C (clk), .D (new_AGEMA_signal_22730), .Q (new_AGEMA_signal_22731) ) ;
    buf_clk new_AGEMA_reg_buffer_10011 ( .C (clk), .D (new_AGEMA_signal_22734), .Q (new_AGEMA_signal_22735) ) ;
    buf_clk new_AGEMA_reg_buffer_10015 ( .C (clk), .D (new_AGEMA_signal_22738), .Q (new_AGEMA_signal_22739) ) ;
    buf_clk new_AGEMA_reg_buffer_10019 ( .C (clk), .D (new_AGEMA_signal_22742), .Q (new_AGEMA_signal_22743) ) ;
    buf_clk new_AGEMA_reg_buffer_10023 ( .C (clk), .D (new_AGEMA_signal_22746), .Q (new_AGEMA_signal_22747) ) ;
    buf_clk new_AGEMA_reg_buffer_10027 ( .C (clk), .D (new_AGEMA_signal_22750), .Q (new_AGEMA_signal_22751) ) ;
    buf_clk new_AGEMA_reg_buffer_10031 ( .C (clk), .D (new_AGEMA_signal_22754), .Q (new_AGEMA_signal_22755) ) ;
    buf_clk new_AGEMA_reg_buffer_10035 ( .C (clk), .D (new_AGEMA_signal_22758), .Q (new_AGEMA_signal_22759) ) ;
    buf_clk new_AGEMA_reg_buffer_10039 ( .C (clk), .D (new_AGEMA_signal_22762), .Q (new_AGEMA_signal_22763) ) ;
    buf_clk new_AGEMA_reg_buffer_10043 ( .C (clk), .D (new_AGEMA_signal_22766), .Q (new_AGEMA_signal_22767) ) ;
    buf_clk new_AGEMA_reg_buffer_10047 ( .C (clk), .D (new_AGEMA_signal_22770), .Q (new_AGEMA_signal_22771) ) ;
    buf_clk new_AGEMA_reg_buffer_10051 ( .C (clk), .D (new_AGEMA_signal_22774), .Q (new_AGEMA_signal_22775) ) ;
    buf_clk new_AGEMA_reg_buffer_10055 ( .C (clk), .D (new_AGEMA_signal_22778), .Q (new_AGEMA_signal_22779) ) ;
    buf_clk new_AGEMA_reg_buffer_10059 ( .C (clk), .D (new_AGEMA_signal_22782), .Q (new_AGEMA_signal_22783) ) ;
    buf_clk new_AGEMA_reg_buffer_10063 ( .C (clk), .D (new_AGEMA_signal_22786), .Q (new_AGEMA_signal_22787) ) ;
    buf_clk new_AGEMA_reg_buffer_10067 ( .C (clk), .D (new_AGEMA_signal_22790), .Q (new_AGEMA_signal_22791) ) ;
    buf_clk new_AGEMA_reg_buffer_10071 ( .C (clk), .D (new_AGEMA_signal_22794), .Q (new_AGEMA_signal_22795) ) ;
    buf_clk new_AGEMA_reg_buffer_10075 ( .C (clk), .D (new_AGEMA_signal_22798), .Q (new_AGEMA_signal_22799) ) ;
    buf_clk new_AGEMA_reg_buffer_10079 ( .C (clk), .D (new_AGEMA_signal_22802), .Q (new_AGEMA_signal_22803) ) ;
    buf_clk new_AGEMA_reg_buffer_10083 ( .C (clk), .D (new_AGEMA_signal_22806), .Q (new_AGEMA_signal_22807) ) ;
    buf_clk new_AGEMA_reg_buffer_10087 ( .C (clk), .D (new_AGEMA_signal_22810), .Q (new_AGEMA_signal_22811) ) ;
    buf_clk new_AGEMA_reg_buffer_10091 ( .C (clk), .D (new_AGEMA_signal_22814), .Q (new_AGEMA_signal_22815) ) ;
    buf_clk new_AGEMA_reg_buffer_10095 ( .C (clk), .D (new_AGEMA_signal_22818), .Q (new_AGEMA_signal_22819) ) ;
    buf_clk new_AGEMA_reg_buffer_10099 ( .C (clk), .D (new_AGEMA_signal_22822), .Q (new_AGEMA_signal_22823) ) ;
    buf_clk new_AGEMA_reg_buffer_10103 ( .C (clk), .D (new_AGEMA_signal_22826), .Q (new_AGEMA_signal_22827) ) ;
    buf_clk new_AGEMA_reg_buffer_10107 ( .C (clk), .D (new_AGEMA_signal_22830), .Q (new_AGEMA_signal_22831) ) ;
    buf_clk new_AGEMA_reg_buffer_10111 ( .C (clk), .D (new_AGEMA_signal_22834), .Q (new_AGEMA_signal_22835) ) ;
    buf_clk new_AGEMA_reg_buffer_10115 ( .C (clk), .D (new_AGEMA_signal_22838), .Q (new_AGEMA_signal_22839) ) ;
    buf_clk new_AGEMA_reg_buffer_10119 ( .C (clk), .D (new_AGEMA_signal_22842), .Q (new_AGEMA_signal_22843) ) ;
    buf_clk new_AGEMA_reg_buffer_10123 ( .C (clk), .D (new_AGEMA_signal_22846), .Q (new_AGEMA_signal_22847) ) ;
    buf_clk new_AGEMA_reg_buffer_10127 ( .C (clk), .D (new_AGEMA_signal_22850), .Q (new_AGEMA_signal_22851) ) ;
    buf_clk new_AGEMA_reg_buffer_10131 ( .C (clk), .D (new_AGEMA_signal_22854), .Q (new_AGEMA_signal_22855) ) ;
    buf_clk new_AGEMA_reg_buffer_10135 ( .C (clk), .D (new_AGEMA_signal_22858), .Q (new_AGEMA_signal_22859) ) ;
    buf_clk new_AGEMA_reg_buffer_10139 ( .C (clk), .D (new_AGEMA_signal_22862), .Q (new_AGEMA_signal_22863) ) ;
    buf_clk new_AGEMA_reg_buffer_10143 ( .C (clk), .D (new_AGEMA_signal_22866), .Q (new_AGEMA_signal_22867) ) ;
    buf_clk new_AGEMA_reg_buffer_10147 ( .C (clk), .D (new_AGEMA_signal_22870), .Q (new_AGEMA_signal_22871) ) ;
    buf_clk new_AGEMA_reg_buffer_10151 ( .C (clk), .D (new_AGEMA_signal_22874), .Q (new_AGEMA_signal_22875) ) ;
    buf_clk new_AGEMA_reg_buffer_10155 ( .C (clk), .D (new_AGEMA_signal_22878), .Q (new_AGEMA_signal_22879) ) ;
    buf_clk new_AGEMA_reg_buffer_10159 ( .C (clk), .D (new_AGEMA_signal_22882), .Q (new_AGEMA_signal_22883) ) ;
    buf_clk new_AGEMA_reg_buffer_10163 ( .C (clk), .D (new_AGEMA_signal_22886), .Q (new_AGEMA_signal_22887) ) ;
    buf_clk new_AGEMA_reg_buffer_10167 ( .C (clk), .D (new_AGEMA_signal_22890), .Q (new_AGEMA_signal_22891) ) ;
    buf_clk new_AGEMA_reg_buffer_10171 ( .C (clk), .D (new_AGEMA_signal_22894), .Q (new_AGEMA_signal_22895) ) ;
    buf_clk new_AGEMA_reg_buffer_10175 ( .C (clk), .D (new_AGEMA_signal_22898), .Q (new_AGEMA_signal_22899) ) ;
    buf_clk new_AGEMA_reg_buffer_10179 ( .C (clk), .D (new_AGEMA_signal_22902), .Q (new_AGEMA_signal_22903) ) ;
    buf_clk new_AGEMA_reg_buffer_10183 ( .C (clk), .D (new_AGEMA_signal_22906), .Q (new_AGEMA_signal_22907) ) ;
    buf_clk new_AGEMA_reg_buffer_10187 ( .C (clk), .D (new_AGEMA_signal_22910), .Q (new_AGEMA_signal_22911) ) ;
    buf_clk new_AGEMA_reg_buffer_10191 ( .C (clk), .D (new_AGEMA_signal_22914), .Q (new_AGEMA_signal_22915) ) ;
    buf_clk new_AGEMA_reg_buffer_10195 ( .C (clk), .D (new_AGEMA_signal_22918), .Q (new_AGEMA_signal_22919) ) ;
    buf_clk new_AGEMA_reg_buffer_10199 ( .C (clk), .D (new_AGEMA_signal_22922), .Q (new_AGEMA_signal_22923) ) ;
    buf_clk new_AGEMA_reg_buffer_10203 ( .C (clk), .D (new_AGEMA_signal_22926), .Q (new_AGEMA_signal_22927) ) ;
    buf_clk new_AGEMA_reg_buffer_10207 ( .C (clk), .D (new_AGEMA_signal_22930), .Q (new_AGEMA_signal_22931) ) ;
    buf_clk new_AGEMA_reg_buffer_10211 ( .C (clk), .D (new_AGEMA_signal_22934), .Q (new_AGEMA_signal_22935) ) ;
    buf_clk new_AGEMA_reg_buffer_10215 ( .C (clk), .D (new_AGEMA_signal_22938), .Q (new_AGEMA_signal_22939) ) ;
    buf_clk new_AGEMA_reg_buffer_10219 ( .C (clk), .D (new_AGEMA_signal_22942), .Q (new_AGEMA_signal_22943) ) ;
    buf_clk new_AGEMA_reg_buffer_10223 ( .C (clk), .D (new_AGEMA_signal_22946), .Q (new_AGEMA_signal_22947) ) ;
    buf_clk new_AGEMA_reg_buffer_10227 ( .C (clk), .D (new_AGEMA_signal_22950), .Q (new_AGEMA_signal_22951) ) ;
    buf_clk new_AGEMA_reg_buffer_10231 ( .C (clk), .D (new_AGEMA_signal_22954), .Q (new_AGEMA_signal_22955) ) ;
    buf_clk new_AGEMA_reg_buffer_10235 ( .C (clk), .D (new_AGEMA_signal_22958), .Q (new_AGEMA_signal_22959) ) ;
    buf_clk new_AGEMA_reg_buffer_10239 ( .C (clk), .D (new_AGEMA_signal_22962), .Q (new_AGEMA_signal_22963) ) ;
    buf_clk new_AGEMA_reg_buffer_10243 ( .C (clk), .D (new_AGEMA_signal_22966), .Q (new_AGEMA_signal_22967) ) ;
    buf_clk new_AGEMA_reg_buffer_10247 ( .C (clk), .D (new_AGEMA_signal_22970), .Q (new_AGEMA_signal_22971) ) ;
    buf_clk new_AGEMA_reg_buffer_10251 ( .C (clk), .D (new_AGEMA_signal_22974), .Q (new_AGEMA_signal_22975) ) ;
    buf_clk new_AGEMA_reg_buffer_10255 ( .C (clk), .D (new_AGEMA_signal_22978), .Q (new_AGEMA_signal_22979) ) ;
    buf_clk new_AGEMA_reg_buffer_10259 ( .C (clk), .D (new_AGEMA_signal_22982), .Q (new_AGEMA_signal_22983) ) ;
    buf_clk new_AGEMA_reg_buffer_10263 ( .C (clk), .D (new_AGEMA_signal_22986), .Q (new_AGEMA_signal_22987) ) ;
    buf_clk new_AGEMA_reg_buffer_10267 ( .C (clk), .D (new_AGEMA_signal_22990), .Q (new_AGEMA_signal_22991) ) ;
    buf_clk new_AGEMA_reg_buffer_10271 ( .C (clk), .D (new_AGEMA_signal_22994), .Q (new_AGEMA_signal_22995) ) ;
    buf_clk new_AGEMA_reg_buffer_10275 ( .C (clk), .D (new_AGEMA_signal_22998), .Q (new_AGEMA_signal_22999) ) ;
    buf_clk new_AGEMA_reg_buffer_10279 ( .C (clk), .D (new_AGEMA_signal_23002), .Q (new_AGEMA_signal_23003) ) ;
    buf_clk new_AGEMA_reg_buffer_10283 ( .C (clk), .D (new_AGEMA_signal_23006), .Q (new_AGEMA_signal_23007) ) ;
    buf_clk new_AGEMA_reg_buffer_10287 ( .C (clk), .D (new_AGEMA_signal_23010), .Q (new_AGEMA_signal_23011) ) ;
    buf_clk new_AGEMA_reg_buffer_10291 ( .C (clk), .D (new_AGEMA_signal_23014), .Q (new_AGEMA_signal_23015) ) ;
    buf_clk new_AGEMA_reg_buffer_10295 ( .C (clk), .D (new_AGEMA_signal_23018), .Q (new_AGEMA_signal_23019) ) ;
    buf_clk new_AGEMA_reg_buffer_10299 ( .C (clk), .D (new_AGEMA_signal_23022), .Q (new_AGEMA_signal_23023) ) ;
    buf_clk new_AGEMA_reg_buffer_10303 ( .C (clk), .D (new_AGEMA_signal_23026), .Q (new_AGEMA_signal_23027) ) ;
    buf_clk new_AGEMA_reg_buffer_10307 ( .C (clk), .D (new_AGEMA_signal_23030), .Q (new_AGEMA_signal_23031) ) ;
    buf_clk new_AGEMA_reg_buffer_10311 ( .C (clk), .D (new_AGEMA_signal_23034), .Q (new_AGEMA_signal_23035) ) ;
    buf_clk new_AGEMA_reg_buffer_10315 ( .C (clk), .D (new_AGEMA_signal_23038), .Q (new_AGEMA_signal_23039) ) ;
    buf_clk new_AGEMA_reg_buffer_10319 ( .C (clk), .D (new_AGEMA_signal_23042), .Q (new_AGEMA_signal_23043) ) ;
    buf_clk new_AGEMA_reg_buffer_10323 ( .C (clk), .D (new_AGEMA_signal_23046), .Q (new_AGEMA_signal_23047) ) ;
    buf_clk new_AGEMA_reg_buffer_10327 ( .C (clk), .D (new_AGEMA_signal_23050), .Q (new_AGEMA_signal_23051) ) ;
    buf_clk new_AGEMA_reg_buffer_10331 ( .C (clk), .D (new_AGEMA_signal_23054), .Q (new_AGEMA_signal_23055) ) ;
    buf_clk new_AGEMA_reg_buffer_10335 ( .C (clk), .D (new_AGEMA_signal_23058), .Q (new_AGEMA_signal_23059) ) ;
    buf_clk new_AGEMA_reg_buffer_10339 ( .C (clk), .D (new_AGEMA_signal_23062), .Q (new_AGEMA_signal_23063) ) ;
    buf_clk new_AGEMA_reg_buffer_10343 ( .C (clk), .D (new_AGEMA_signal_23066), .Q (new_AGEMA_signal_23067) ) ;
    buf_clk new_AGEMA_reg_buffer_10347 ( .C (clk), .D (new_AGEMA_signal_23070), .Q (new_AGEMA_signal_23071) ) ;
    buf_clk new_AGEMA_reg_buffer_10351 ( .C (clk), .D (new_AGEMA_signal_23074), .Q (new_AGEMA_signal_23075) ) ;
    buf_clk new_AGEMA_reg_buffer_10355 ( .C (clk), .D (new_AGEMA_signal_23078), .Q (new_AGEMA_signal_23079) ) ;
    buf_clk new_AGEMA_reg_buffer_10359 ( .C (clk), .D (new_AGEMA_signal_23082), .Q (new_AGEMA_signal_23083) ) ;
    buf_clk new_AGEMA_reg_buffer_10363 ( .C (clk), .D (new_AGEMA_signal_23086), .Q (new_AGEMA_signal_23087) ) ;
    buf_clk new_AGEMA_reg_buffer_10367 ( .C (clk), .D (new_AGEMA_signal_23090), .Q (new_AGEMA_signal_23091) ) ;
    buf_clk new_AGEMA_reg_buffer_10371 ( .C (clk), .D (new_AGEMA_signal_23094), .Q (new_AGEMA_signal_23095) ) ;
    buf_clk new_AGEMA_reg_buffer_10375 ( .C (clk), .D (new_AGEMA_signal_23098), .Q (new_AGEMA_signal_23099) ) ;
    buf_clk new_AGEMA_reg_buffer_10379 ( .C (clk), .D (new_AGEMA_signal_23102), .Q (new_AGEMA_signal_23103) ) ;
    buf_clk new_AGEMA_reg_buffer_10383 ( .C (clk), .D (new_AGEMA_signal_23106), .Q (new_AGEMA_signal_23107) ) ;
    buf_clk new_AGEMA_reg_buffer_10387 ( .C (clk), .D (new_AGEMA_signal_23110), .Q (new_AGEMA_signal_23111) ) ;
    buf_clk new_AGEMA_reg_buffer_10391 ( .C (clk), .D (new_AGEMA_signal_23114), .Q (new_AGEMA_signal_23115) ) ;
    buf_clk new_AGEMA_reg_buffer_10395 ( .C (clk), .D (new_AGEMA_signal_23118), .Q (new_AGEMA_signal_23119) ) ;
    buf_clk new_AGEMA_reg_buffer_10399 ( .C (clk), .D (new_AGEMA_signal_23122), .Q (new_AGEMA_signal_23123) ) ;
    buf_clk new_AGEMA_reg_buffer_10403 ( .C (clk), .D (new_AGEMA_signal_23126), .Q (new_AGEMA_signal_23127) ) ;
    buf_clk new_AGEMA_reg_buffer_10407 ( .C (clk), .D (new_AGEMA_signal_23130), .Q (new_AGEMA_signal_23131) ) ;
    buf_clk new_AGEMA_reg_buffer_10411 ( .C (clk), .D (new_AGEMA_signal_23134), .Q (new_AGEMA_signal_23135) ) ;
    buf_clk new_AGEMA_reg_buffer_10415 ( .C (clk), .D (new_AGEMA_signal_23138), .Q (new_AGEMA_signal_23139) ) ;
    buf_clk new_AGEMA_reg_buffer_10419 ( .C (clk), .D (new_AGEMA_signal_23142), .Q (new_AGEMA_signal_23143) ) ;
    buf_clk new_AGEMA_reg_buffer_10423 ( .C (clk), .D (new_AGEMA_signal_23146), .Q (new_AGEMA_signal_23147) ) ;
    buf_clk new_AGEMA_reg_buffer_10427 ( .C (clk), .D (new_AGEMA_signal_23150), .Q (new_AGEMA_signal_23151) ) ;
    buf_clk new_AGEMA_reg_buffer_10431 ( .C (clk), .D (new_AGEMA_signal_23154), .Q (new_AGEMA_signal_23155) ) ;
    buf_clk new_AGEMA_reg_buffer_10435 ( .C (clk), .D (new_AGEMA_signal_23158), .Q (new_AGEMA_signal_23159) ) ;
    buf_clk new_AGEMA_reg_buffer_10439 ( .C (clk), .D (new_AGEMA_signal_23162), .Q (new_AGEMA_signal_23163) ) ;
    buf_clk new_AGEMA_reg_buffer_10443 ( .C (clk), .D (new_AGEMA_signal_23166), .Q (new_AGEMA_signal_23167) ) ;
    buf_clk new_AGEMA_reg_buffer_10447 ( .C (clk), .D (new_AGEMA_signal_23170), .Q (new_AGEMA_signal_23171) ) ;
    buf_clk new_AGEMA_reg_buffer_10451 ( .C (clk), .D (new_AGEMA_signal_23174), .Q (new_AGEMA_signal_23175) ) ;
    buf_clk new_AGEMA_reg_buffer_10455 ( .C (clk), .D (new_AGEMA_signal_23178), .Q (new_AGEMA_signal_23179) ) ;
    buf_clk new_AGEMA_reg_buffer_10459 ( .C (clk), .D (new_AGEMA_signal_23182), .Q (new_AGEMA_signal_23183) ) ;
    buf_clk new_AGEMA_reg_buffer_10463 ( .C (clk), .D (new_AGEMA_signal_23186), .Q (new_AGEMA_signal_23187) ) ;
    buf_clk new_AGEMA_reg_buffer_10467 ( .C (clk), .D (new_AGEMA_signal_23190), .Q (new_AGEMA_signal_23191) ) ;
    buf_clk new_AGEMA_reg_buffer_10471 ( .C (clk), .D (new_AGEMA_signal_23194), .Q (new_AGEMA_signal_23195) ) ;
    buf_clk new_AGEMA_reg_buffer_10475 ( .C (clk), .D (new_AGEMA_signal_23198), .Q (new_AGEMA_signal_23199) ) ;
    buf_clk new_AGEMA_reg_buffer_10479 ( .C (clk), .D (new_AGEMA_signal_23202), .Q (new_AGEMA_signal_23203) ) ;
    buf_clk new_AGEMA_reg_buffer_10483 ( .C (clk), .D (new_AGEMA_signal_23206), .Q (new_AGEMA_signal_23207) ) ;
    buf_clk new_AGEMA_reg_buffer_10487 ( .C (clk), .D (new_AGEMA_signal_23210), .Q (new_AGEMA_signal_23211) ) ;
    buf_clk new_AGEMA_reg_buffer_10491 ( .C (clk), .D (new_AGEMA_signal_23214), .Q (new_AGEMA_signal_23215) ) ;
    buf_clk new_AGEMA_reg_buffer_10495 ( .C (clk), .D (new_AGEMA_signal_23218), .Q (new_AGEMA_signal_23219) ) ;
    buf_clk new_AGEMA_reg_buffer_10499 ( .C (clk), .D (new_AGEMA_signal_23222), .Q (new_AGEMA_signal_23223) ) ;
    buf_clk new_AGEMA_reg_buffer_10503 ( .C (clk), .D (new_AGEMA_signal_23226), .Q (new_AGEMA_signal_23227) ) ;
    buf_clk new_AGEMA_reg_buffer_10507 ( .C (clk), .D (new_AGEMA_signal_23230), .Q (new_AGEMA_signal_23231) ) ;
    buf_clk new_AGEMA_reg_buffer_10511 ( .C (clk), .D (new_AGEMA_signal_23234), .Q (new_AGEMA_signal_23235) ) ;
    buf_clk new_AGEMA_reg_buffer_10515 ( .C (clk), .D (new_AGEMA_signal_23238), .Q (new_AGEMA_signal_23239) ) ;
    buf_clk new_AGEMA_reg_buffer_10519 ( .C (clk), .D (new_AGEMA_signal_23242), .Q (new_AGEMA_signal_23243) ) ;
    buf_clk new_AGEMA_reg_buffer_10523 ( .C (clk), .D (new_AGEMA_signal_23246), .Q (new_AGEMA_signal_23247) ) ;
    buf_clk new_AGEMA_reg_buffer_10527 ( .C (clk), .D (new_AGEMA_signal_23250), .Q (new_AGEMA_signal_23251) ) ;
    buf_clk new_AGEMA_reg_buffer_10531 ( .C (clk), .D (new_AGEMA_signal_23254), .Q (new_AGEMA_signal_23255) ) ;
    buf_clk new_AGEMA_reg_buffer_10535 ( .C (clk), .D (new_AGEMA_signal_23258), .Q (new_AGEMA_signal_23259) ) ;
    buf_clk new_AGEMA_reg_buffer_10539 ( .C (clk), .D (new_AGEMA_signal_23262), .Q (new_AGEMA_signal_23263) ) ;
    buf_clk new_AGEMA_reg_buffer_10543 ( .C (clk), .D (new_AGEMA_signal_23266), .Q (new_AGEMA_signal_23267) ) ;
    buf_clk new_AGEMA_reg_buffer_10547 ( .C (clk), .D (new_AGEMA_signal_23270), .Q (new_AGEMA_signal_23271) ) ;
    buf_clk new_AGEMA_reg_buffer_10551 ( .C (clk), .D (new_AGEMA_signal_23274), .Q (new_AGEMA_signal_23275) ) ;
    buf_clk new_AGEMA_reg_buffer_10555 ( .C (clk), .D (new_AGEMA_signal_23278), .Q (new_AGEMA_signal_23279) ) ;
    buf_clk new_AGEMA_reg_buffer_10559 ( .C (clk), .D (new_AGEMA_signal_23282), .Q (new_AGEMA_signal_23283) ) ;
    buf_clk new_AGEMA_reg_buffer_10563 ( .C (clk), .D (new_AGEMA_signal_23286), .Q (new_AGEMA_signal_23287) ) ;
    buf_clk new_AGEMA_reg_buffer_10567 ( .C (clk), .D (new_AGEMA_signal_23290), .Q (new_AGEMA_signal_23291) ) ;
    buf_clk new_AGEMA_reg_buffer_10571 ( .C (clk), .D (new_AGEMA_signal_23294), .Q (new_AGEMA_signal_23295) ) ;
    buf_clk new_AGEMA_reg_buffer_10575 ( .C (clk), .D (new_AGEMA_signal_23298), .Q (new_AGEMA_signal_23299) ) ;
    buf_clk new_AGEMA_reg_buffer_10579 ( .C (clk), .D (new_AGEMA_signal_23302), .Q (new_AGEMA_signal_23303) ) ;
    buf_clk new_AGEMA_reg_buffer_10583 ( .C (clk), .D (new_AGEMA_signal_23306), .Q (new_AGEMA_signal_23307) ) ;
    buf_clk new_AGEMA_reg_buffer_10587 ( .C (clk), .D (new_AGEMA_signal_23310), .Q (new_AGEMA_signal_23311) ) ;
    buf_clk new_AGEMA_reg_buffer_10591 ( .C (clk), .D (new_AGEMA_signal_23314), .Q (new_AGEMA_signal_23315) ) ;
    buf_clk new_AGEMA_reg_buffer_10595 ( .C (clk), .D (new_AGEMA_signal_23318), .Q (new_AGEMA_signal_23319) ) ;
    buf_clk new_AGEMA_reg_buffer_10599 ( .C (clk), .D (new_AGEMA_signal_23322), .Q (new_AGEMA_signal_23323) ) ;
    buf_clk new_AGEMA_reg_buffer_10603 ( .C (clk), .D (new_AGEMA_signal_23326), .Q (new_AGEMA_signal_23327) ) ;
    buf_clk new_AGEMA_reg_buffer_10607 ( .C (clk), .D (new_AGEMA_signal_23330), .Q (new_AGEMA_signal_23331) ) ;
    buf_clk new_AGEMA_reg_buffer_10611 ( .C (clk), .D (new_AGEMA_signal_23334), .Q (new_AGEMA_signal_23335) ) ;
    buf_clk new_AGEMA_reg_buffer_10615 ( .C (clk), .D (new_AGEMA_signal_23338), .Q (new_AGEMA_signal_23339) ) ;
    buf_clk new_AGEMA_reg_buffer_10619 ( .C (clk), .D (new_AGEMA_signal_23342), .Q (new_AGEMA_signal_23343) ) ;
    buf_clk new_AGEMA_reg_buffer_10623 ( .C (clk), .D (new_AGEMA_signal_23346), .Q (new_AGEMA_signal_23347) ) ;
    buf_clk new_AGEMA_reg_buffer_10627 ( .C (clk), .D (new_AGEMA_signal_23350), .Q (new_AGEMA_signal_23351) ) ;
    buf_clk new_AGEMA_reg_buffer_10631 ( .C (clk), .D (new_AGEMA_signal_23354), .Q (new_AGEMA_signal_23355) ) ;
    buf_clk new_AGEMA_reg_buffer_10635 ( .C (clk), .D (new_AGEMA_signal_23358), .Q (new_AGEMA_signal_23359) ) ;
    buf_clk new_AGEMA_reg_buffer_10639 ( .C (clk), .D (new_AGEMA_signal_23362), .Q (new_AGEMA_signal_23363) ) ;
    buf_clk new_AGEMA_reg_buffer_10643 ( .C (clk), .D (new_AGEMA_signal_23366), .Q (new_AGEMA_signal_23367) ) ;
    buf_clk new_AGEMA_reg_buffer_10647 ( .C (clk), .D (new_AGEMA_signal_23370), .Q (new_AGEMA_signal_23371) ) ;
    buf_clk new_AGEMA_reg_buffer_10651 ( .C (clk), .D (new_AGEMA_signal_23374), .Q (new_AGEMA_signal_23375) ) ;
    buf_clk new_AGEMA_reg_buffer_10655 ( .C (clk), .D (new_AGEMA_signal_23378), .Q (new_AGEMA_signal_23379) ) ;
    buf_clk new_AGEMA_reg_buffer_10659 ( .C (clk), .D (new_AGEMA_signal_23382), .Q (new_AGEMA_signal_23383) ) ;
    buf_clk new_AGEMA_reg_buffer_10663 ( .C (clk), .D (new_AGEMA_signal_23386), .Q (new_AGEMA_signal_23387) ) ;
    buf_clk new_AGEMA_reg_buffer_10667 ( .C (clk), .D (new_AGEMA_signal_23390), .Q (new_AGEMA_signal_23391) ) ;
    buf_clk new_AGEMA_reg_buffer_10671 ( .C (clk), .D (new_AGEMA_signal_23394), .Q (new_AGEMA_signal_23395) ) ;
    buf_clk new_AGEMA_reg_buffer_10675 ( .C (clk), .D (new_AGEMA_signal_23398), .Q (new_AGEMA_signal_23399) ) ;
    buf_clk new_AGEMA_reg_buffer_10679 ( .C (clk), .D (new_AGEMA_signal_23402), .Q (new_AGEMA_signal_23403) ) ;
    buf_clk new_AGEMA_reg_buffer_10683 ( .C (clk), .D (new_AGEMA_signal_23406), .Q (new_AGEMA_signal_23407) ) ;
    buf_clk new_AGEMA_reg_buffer_10687 ( .C (clk), .D (new_AGEMA_signal_23410), .Q (new_AGEMA_signal_23411) ) ;
    buf_clk new_AGEMA_reg_buffer_10691 ( .C (clk), .D (new_AGEMA_signal_23414), .Q (new_AGEMA_signal_23415) ) ;
    buf_clk new_AGEMA_reg_buffer_10695 ( .C (clk), .D (new_AGEMA_signal_23418), .Q (new_AGEMA_signal_23419) ) ;
    buf_clk new_AGEMA_reg_buffer_10699 ( .C (clk), .D (new_AGEMA_signal_23422), .Q (new_AGEMA_signal_23423) ) ;
    buf_clk new_AGEMA_reg_buffer_10703 ( .C (clk), .D (new_AGEMA_signal_23426), .Q (new_AGEMA_signal_23427) ) ;
    buf_clk new_AGEMA_reg_buffer_10707 ( .C (clk), .D (new_AGEMA_signal_23430), .Q (new_AGEMA_signal_23431) ) ;
    buf_clk new_AGEMA_reg_buffer_10711 ( .C (clk), .D (new_AGEMA_signal_23434), .Q (new_AGEMA_signal_23435) ) ;
    buf_clk new_AGEMA_reg_buffer_10715 ( .C (clk), .D (new_AGEMA_signal_23438), .Q (new_AGEMA_signal_23439) ) ;
    buf_clk new_AGEMA_reg_buffer_10719 ( .C (clk), .D (new_AGEMA_signal_23442), .Q (new_AGEMA_signal_23443) ) ;
    buf_clk new_AGEMA_reg_buffer_10723 ( .C (clk), .D (new_AGEMA_signal_23446), .Q (new_AGEMA_signal_23447) ) ;
    buf_clk new_AGEMA_reg_buffer_10727 ( .C (clk), .D (new_AGEMA_signal_23450), .Q (new_AGEMA_signal_23451) ) ;
    buf_clk new_AGEMA_reg_buffer_10731 ( .C (clk), .D (new_AGEMA_signal_23454), .Q (new_AGEMA_signal_23455) ) ;
    buf_clk new_AGEMA_reg_buffer_10735 ( .C (clk), .D (new_AGEMA_signal_23458), .Q (new_AGEMA_signal_23459) ) ;
    buf_clk new_AGEMA_reg_buffer_10739 ( .C (clk), .D (new_AGEMA_signal_23462), .Q (new_AGEMA_signal_23463) ) ;
    buf_clk new_AGEMA_reg_buffer_10743 ( .C (clk), .D (new_AGEMA_signal_23466), .Q (new_AGEMA_signal_23467) ) ;
    buf_clk new_AGEMA_reg_buffer_10747 ( .C (clk), .D (new_AGEMA_signal_23470), .Q (new_AGEMA_signal_23471) ) ;
    buf_clk new_AGEMA_reg_buffer_10751 ( .C (clk), .D (new_AGEMA_signal_23474), .Q (new_AGEMA_signal_23475) ) ;
    buf_clk new_AGEMA_reg_buffer_10755 ( .C (clk), .D (new_AGEMA_signal_23478), .Q (new_AGEMA_signal_23479) ) ;
    buf_clk new_AGEMA_reg_buffer_10759 ( .C (clk), .D (new_AGEMA_signal_23482), .Q (new_AGEMA_signal_23483) ) ;
    buf_clk new_AGEMA_reg_buffer_10763 ( .C (clk), .D (new_AGEMA_signal_23486), .Q (new_AGEMA_signal_23487) ) ;
    buf_clk new_AGEMA_reg_buffer_10767 ( .C (clk), .D (new_AGEMA_signal_23490), .Q (new_AGEMA_signal_23491) ) ;
    buf_clk new_AGEMA_reg_buffer_10771 ( .C (clk), .D (new_AGEMA_signal_23494), .Q (new_AGEMA_signal_23495) ) ;
    buf_clk new_AGEMA_reg_buffer_10775 ( .C (clk), .D (new_AGEMA_signal_23498), .Q (new_AGEMA_signal_23499) ) ;
    buf_clk new_AGEMA_reg_buffer_10779 ( .C (clk), .D (new_AGEMA_signal_23502), .Q (new_AGEMA_signal_23503) ) ;
    buf_clk new_AGEMA_reg_buffer_10783 ( .C (clk), .D (new_AGEMA_signal_23506), .Q (new_AGEMA_signal_23507) ) ;
    buf_clk new_AGEMA_reg_buffer_10787 ( .C (clk), .D (new_AGEMA_signal_23510), .Q (new_AGEMA_signal_23511) ) ;
    buf_clk new_AGEMA_reg_buffer_10791 ( .C (clk), .D (new_AGEMA_signal_23514), .Q (new_AGEMA_signal_23515) ) ;
    buf_clk new_AGEMA_reg_buffer_10795 ( .C (clk), .D (new_AGEMA_signal_23518), .Q (new_AGEMA_signal_23519) ) ;
    buf_clk new_AGEMA_reg_buffer_10799 ( .C (clk), .D (new_AGEMA_signal_23522), .Q (new_AGEMA_signal_23523) ) ;
    buf_clk new_AGEMA_reg_buffer_10803 ( .C (clk), .D (new_AGEMA_signal_23526), .Q (new_AGEMA_signal_23527) ) ;
    buf_clk new_AGEMA_reg_buffer_10807 ( .C (clk), .D (new_AGEMA_signal_23530), .Q (new_AGEMA_signal_23531) ) ;
    buf_clk new_AGEMA_reg_buffer_10811 ( .C (clk), .D (new_AGEMA_signal_23534), .Q (new_AGEMA_signal_23535) ) ;
    buf_clk new_AGEMA_reg_buffer_10815 ( .C (clk), .D (new_AGEMA_signal_23538), .Q (new_AGEMA_signal_23539) ) ;
    buf_clk new_AGEMA_reg_buffer_10819 ( .C (clk), .D (new_AGEMA_signal_23542), .Q (new_AGEMA_signal_23543) ) ;
    buf_clk new_AGEMA_reg_buffer_10823 ( .C (clk), .D (new_AGEMA_signal_23546), .Q (new_AGEMA_signal_23547) ) ;
    buf_clk new_AGEMA_reg_buffer_10827 ( .C (clk), .D (new_AGEMA_signal_23550), .Q (new_AGEMA_signal_23551) ) ;
    buf_clk new_AGEMA_reg_buffer_10831 ( .C (clk), .D (new_AGEMA_signal_23554), .Q (new_AGEMA_signal_23555) ) ;
    buf_clk new_AGEMA_reg_buffer_10835 ( .C (clk), .D (new_AGEMA_signal_23558), .Q (new_AGEMA_signal_23559) ) ;
    buf_clk new_AGEMA_reg_buffer_10839 ( .C (clk), .D (new_AGEMA_signal_23562), .Q (new_AGEMA_signal_23563) ) ;
    buf_clk new_AGEMA_reg_buffer_10843 ( .C (clk), .D (new_AGEMA_signal_23566), .Q (new_AGEMA_signal_23567) ) ;
    buf_clk new_AGEMA_reg_buffer_10847 ( .C (clk), .D (new_AGEMA_signal_23570), .Q (new_AGEMA_signal_23571) ) ;
    buf_clk new_AGEMA_reg_buffer_10851 ( .C (clk), .D (new_AGEMA_signal_23574), .Q (new_AGEMA_signal_23575) ) ;
    buf_clk new_AGEMA_reg_buffer_10855 ( .C (clk), .D (new_AGEMA_signal_23578), .Q (new_AGEMA_signal_23579) ) ;
    buf_clk new_AGEMA_reg_buffer_10859 ( .C (clk), .D (new_AGEMA_signal_23582), .Q (new_AGEMA_signal_23583) ) ;
    buf_clk new_AGEMA_reg_buffer_10863 ( .C (clk), .D (new_AGEMA_signal_23586), .Q (new_AGEMA_signal_23587) ) ;
    buf_clk new_AGEMA_reg_buffer_10867 ( .C (clk), .D (new_AGEMA_signal_23590), .Q (new_AGEMA_signal_23591) ) ;
    buf_clk new_AGEMA_reg_buffer_10871 ( .C (clk), .D (new_AGEMA_signal_23594), .Q (new_AGEMA_signal_23595) ) ;
    buf_clk new_AGEMA_reg_buffer_10875 ( .C (clk), .D (new_AGEMA_signal_23598), .Q (new_AGEMA_signal_23599) ) ;
    buf_clk new_AGEMA_reg_buffer_10879 ( .C (clk), .D (new_AGEMA_signal_23602), .Q (new_AGEMA_signal_23603) ) ;
    buf_clk new_AGEMA_reg_buffer_10883 ( .C (clk), .D (new_AGEMA_signal_23606), .Q (new_AGEMA_signal_23607) ) ;
    buf_clk new_AGEMA_reg_buffer_10887 ( .C (clk), .D (new_AGEMA_signal_23610), .Q (new_AGEMA_signal_23611) ) ;
    buf_clk new_AGEMA_reg_buffer_10891 ( .C (clk), .D (new_AGEMA_signal_23614), .Q (new_AGEMA_signal_23615) ) ;
    buf_clk new_AGEMA_reg_buffer_10895 ( .C (clk), .D (new_AGEMA_signal_23618), .Q (new_AGEMA_signal_23619) ) ;
    buf_clk new_AGEMA_reg_buffer_10899 ( .C (clk), .D (new_AGEMA_signal_23622), .Q (new_AGEMA_signal_23623) ) ;
    buf_clk new_AGEMA_reg_buffer_10903 ( .C (clk), .D (new_AGEMA_signal_23626), .Q (new_AGEMA_signal_23627) ) ;
    buf_clk new_AGEMA_reg_buffer_10907 ( .C (clk), .D (new_AGEMA_signal_23630), .Q (new_AGEMA_signal_23631) ) ;
    buf_clk new_AGEMA_reg_buffer_10911 ( .C (clk), .D (new_AGEMA_signal_23634), .Q (new_AGEMA_signal_23635) ) ;
    buf_clk new_AGEMA_reg_buffer_10915 ( .C (clk), .D (new_AGEMA_signal_23638), .Q (new_AGEMA_signal_23639) ) ;
    buf_clk new_AGEMA_reg_buffer_10919 ( .C (clk), .D (new_AGEMA_signal_23642), .Q (new_AGEMA_signal_23643) ) ;
    buf_clk new_AGEMA_reg_buffer_10923 ( .C (clk), .D (new_AGEMA_signal_23646), .Q (new_AGEMA_signal_23647) ) ;
    buf_clk new_AGEMA_reg_buffer_10927 ( .C (clk), .D (new_AGEMA_signal_23650), .Q (new_AGEMA_signal_23651) ) ;
    buf_clk new_AGEMA_reg_buffer_10931 ( .C (clk), .D (new_AGEMA_signal_23654), .Q (new_AGEMA_signal_23655) ) ;
    buf_clk new_AGEMA_reg_buffer_10935 ( .C (clk), .D (new_AGEMA_signal_23658), .Q (new_AGEMA_signal_23659) ) ;
    buf_clk new_AGEMA_reg_buffer_10939 ( .C (clk), .D (new_AGEMA_signal_23662), .Q (new_AGEMA_signal_23663) ) ;
    buf_clk new_AGEMA_reg_buffer_10943 ( .C (clk), .D (new_AGEMA_signal_23666), .Q (new_AGEMA_signal_23667) ) ;
    buf_clk new_AGEMA_reg_buffer_10947 ( .C (clk), .D (new_AGEMA_signal_23670), .Q (new_AGEMA_signal_23671) ) ;
    buf_clk new_AGEMA_reg_buffer_10951 ( .C (clk), .D (new_AGEMA_signal_23674), .Q (new_AGEMA_signal_23675) ) ;
    buf_clk new_AGEMA_reg_buffer_10955 ( .C (clk), .D (new_AGEMA_signal_23678), .Q (new_AGEMA_signal_23679) ) ;
    buf_clk new_AGEMA_reg_buffer_10959 ( .C (clk), .D (new_AGEMA_signal_23682), .Q (new_AGEMA_signal_23683) ) ;
    buf_clk new_AGEMA_reg_buffer_10963 ( .C (clk), .D (new_AGEMA_signal_23686), .Q (new_AGEMA_signal_23687) ) ;
    buf_clk new_AGEMA_reg_buffer_10967 ( .C (clk), .D (new_AGEMA_signal_23690), .Q (new_AGEMA_signal_23691) ) ;
    buf_clk new_AGEMA_reg_buffer_10971 ( .C (clk), .D (new_AGEMA_signal_23694), .Q (new_AGEMA_signal_23695) ) ;
    buf_clk new_AGEMA_reg_buffer_10975 ( .C (clk), .D (new_AGEMA_signal_23698), .Q (new_AGEMA_signal_23699) ) ;
    buf_clk new_AGEMA_reg_buffer_10979 ( .C (clk), .D (new_AGEMA_signal_23702), .Q (new_AGEMA_signal_23703) ) ;
    buf_clk new_AGEMA_reg_buffer_10983 ( .C (clk), .D (new_AGEMA_signal_23706), .Q (new_AGEMA_signal_23707) ) ;
    buf_clk new_AGEMA_reg_buffer_10987 ( .C (clk), .D (new_AGEMA_signal_23710), .Q (new_AGEMA_signal_23711) ) ;
    buf_clk new_AGEMA_reg_buffer_10991 ( .C (clk), .D (new_AGEMA_signal_23714), .Q (new_AGEMA_signal_23715) ) ;
    buf_clk new_AGEMA_reg_buffer_10995 ( .C (clk), .D (new_AGEMA_signal_23718), .Q (new_AGEMA_signal_23719) ) ;
    buf_clk new_AGEMA_reg_buffer_10999 ( .C (clk), .D (new_AGEMA_signal_23722), .Q (new_AGEMA_signal_23723) ) ;
    buf_clk new_AGEMA_reg_buffer_11003 ( .C (clk), .D (new_AGEMA_signal_23726), .Q (new_AGEMA_signal_23727) ) ;
    buf_clk new_AGEMA_reg_buffer_11007 ( .C (clk), .D (new_AGEMA_signal_23730), .Q (new_AGEMA_signal_23731) ) ;
    buf_clk new_AGEMA_reg_buffer_11011 ( .C (clk), .D (new_AGEMA_signal_23734), .Q (new_AGEMA_signal_23735) ) ;
    buf_clk new_AGEMA_reg_buffer_11015 ( .C (clk), .D (new_AGEMA_signal_23738), .Q (new_AGEMA_signal_23739) ) ;
    buf_clk new_AGEMA_reg_buffer_11019 ( .C (clk), .D (new_AGEMA_signal_23742), .Q (new_AGEMA_signal_23743) ) ;
    buf_clk new_AGEMA_reg_buffer_11023 ( .C (clk), .D (new_AGEMA_signal_23746), .Q (new_AGEMA_signal_23747) ) ;
    buf_clk new_AGEMA_reg_buffer_11027 ( .C (clk), .D (new_AGEMA_signal_23750), .Q (new_AGEMA_signal_23751) ) ;
    buf_clk new_AGEMA_reg_buffer_11031 ( .C (clk), .D (new_AGEMA_signal_23754), .Q (new_AGEMA_signal_23755) ) ;
    buf_clk new_AGEMA_reg_buffer_11035 ( .C (clk), .D (new_AGEMA_signal_23758), .Q (new_AGEMA_signal_23759) ) ;
    buf_clk new_AGEMA_reg_buffer_11039 ( .C (clk), .D (new_AGEMA_signal_23762), .Q (new_AGEMA_signal_23763) ) ;
    buf_clk new_AGEMA_reg_buffer_11043 ( .C (clk), .D (new_AGEMA_signal_23766), .Q (new_AGEMA_signal_23767) ) ;
    buf_clk new_AGEMA_reg_buffer_11047 ( .C (clk), .D (new_AGEMA_signal_23770), .Q (new_AGEMA_signal_23771) ) ;
    buf_clk new_AGEMA_reg_buffer_11051 ( .C (clk), .D (new_AGEMA_signal_23774), .Q (new_AGEMA_signal_23775) ) ;
    buf_clk new_AGEMA_reg_buffer_11055 ( .C (clk), .D (new_AGEMA_signal_23778), .Q (new_AGEMA_signal_23779) ) ;
    buf_clk new_AGEMA_reg_buffer_11059 ( .C (clk), .D (new_AGEMA_signal_23782), .Q (new_AGEMA_signal_23783) ) ;
    buf_clk new_AGEMA_reg_buffer_11063 ( .C (clk), .D (new_AGEMA_signal_23786), .Q (new_AGEMA_signal_23787) ) ;
    buf_clk new_AGEMA_reg_buffer_11067 ( .C (clk), .D (new_AGEMA_signal_23790), .Q (new_AGEMA_signal_23791) ) ;
    buf_clk new_AGEMA_reg_buffer_11071 ( .C (clk), .D (new_AGEMA_signal_23794), .Q (new_AGEMA_signal_23795) ) ;
    buf_clk new_AGEMA_reg_buffer_11075 ( .C (clk), .D (new_AGEMA_signal_23798), .Q (new_AGEMA_signal_23799) ) ;
    buf_clk new_AGEMA_reg_buffer_11079 ( .C (clk), .D (new_AGEMA_signal_23802), .Q (new_AGEMA_signal_23803) ) ;
    buf_clk new_AGEMA_reg_buffer_11083 ( .C (clk), .D (new_AGEMA_signal_23806), .Q (new_AGEMA_signal_23807) ) ;
    buf_clk new_AGEMA_reg_buffer_11087 ( .C (clk), .D (new_AGEMA_signal_23810), .Q (new_AGEMA_signal_23811) ) ;
    buf_clk new_AGEMA_reg_buffer_11091 ( .C (clk), .D (new_AGEMA_signal_23814), .Q (new_AGEMA_signal_23815) ) ;
    buf_clk new_AGEMA_reg_buffer_11095 ( .C (clk), .D (new_AGEMA_signal_23818), .Q (new_AGEMA_signal_23819) ) ;
    buf_clk new_AGEMA_reg_buffer_11099 ( .C (clk), .D (new_AGEMA_signal_23822), .Q (new_AGEMA_signal_23823) ) ;
    buf_clk new_AGEMA_reg_buffer_11103 ( .C (clk), .D (new_AGEMA_signal_23826), .Q (new_AGEMA_signal_23827) ) ;
    buf_clk new_AGEMA_reg_buffer_11107 ( .C (clk), .D (new_AGEMA_signal_23830), .Q (new_AGEMA_signal_23831) ) ;
    buf_clk new_AGEMA_reg_buffer_11111 ( .C (clk), .D (new_AGEMA_signal_23834), .Q (new_AGEMA_signal_23835) ) ;
    buf_clk new_AGEMA_reg_buffer_11115 ( .C (clk), .D (new_AGEMA_signal_23838), .Q (new_AGEMA_signal_23839) ) ;
    buf_clk new_AGEMA_reg_buffer_11119 ( .C (clk), .D (new_AGEMA_signal_23842), .Q (new_AGEMA_signal_23843) ) ;
    buf_clk new_AGEMA_reg_buffer_11123 ( .C (clk), .D (new_AGEMA_signal_23846), .Q (new_AGEMA_signal_23847) ) ;
    buf_clk new_AGEMA_reg_buffer_11127 ( .C (clk), .D (new_AGEMA_signal_23850), .Q (new_AGEMA_signal_23851) ) ;
    buf_clk new_AGEMA_reg_buffer_11131 ( .C (clk), .D (new_AGEMA_signal_23854), .Q (new_AGEMA_signal_23855) ) ;
    buf_clk new_AGEMA_reg_buffer_11135 ( .C (clk), .D (new_AGEMA_signal_23858), .Q (new_AGEMA_signal_23859) ) ;
    buf_clk new_AGEMA_reg_buffer_11139 ( .C (clk), .D (new_AGEMA_signal_23862), .Q (new_AGEMA_signal_23863) ) ;
    buf_clk new_AGEMA_reg_buffer_11143 ( .C (clk), .D (new_AGEMA_signal_23866), .Q (new_AGEMA_signal_23867) ) ;
    buf_clk new_AGEMA_reg_buffer_11147 ( .C (clk), .D (new_AGEMA_signal_23870), .Q (new_AGEMA_signal_23871) ) ;
    buf_clk new_AGEMA_reg_buffer_11151 ( .C (clk), .D (new_AGEMA_signal_23874), .Q (new_AGEMA_signal_23875) ) ;
    buf_clk new_AGEMA_reg_buffer_11155 ( .C (clk), .D (new_AGEMA_signal_23878), .Q (new_AGEMA_signal_23879) ) ;
    buf_clk new_AGEMA_reg_buffer_11159 ( .C (clk), .D (new_AGEMA_signal_23882), .Q (new_AGEMA_signal_23883) ) ;
    buf_clk new_AGEMA_reg_buffer_11163 ( .C (clk), .D (new_AGEMA_signal_23886), .Q (new_AGEMA_signal_23887) ) ;
    buf_clk new_AGEMA_reg_buffer_11167 ( .C (clk), .D (new_AGEMA_signal_23890), .Q (new_AGEMA_signal_23891) ) ;
    buf_clk new_AGEMA_reg_buffer_11171 ( .C (clk), .D (new_AGEMA_signal_23894), .Q (new_AGEMA_signal_23895) ) ;
    buf_clk new_AGEMA_reg_buffer_11175 ( .C (clk), .D (new_AGEMA_signal_23898), .Q (new_AGEMA_signal_23899) ) ;
    buf_clk new_AGEMA_reg_buffer_11179 ( .C (clk), .D (new_AGEMA_signal_23902), .Q (new_AGEMA_signal_23903) ) ;
    buf_clk new_AGEMA_reg_buffer_11183 ( .C (clk), .D (new_AGEMA_signal_23906), .Q (new_AGEMA_signal_23907) ) ;
    buf_clk new_AGEMA_reg_buffer_11187 ( .C (clk), .D (new_AGEMA_signal_23910), .Q (new_AGEMA_signal_23911) ) ;
    buf_clk new_AGEMA_reg_buffer_11191 ( .C (clk), .D (new_AGEMA_signal_23914), .Q (new_AGEMA_signal_23915) ) ;
    buf_clk new_AGEMA_reg_buffer_11195 ( .C (clk), .D (new_AGEMA_signal_23918), .Q (new_AGEMA_signal_23919) ) ;
    buf_clk new_AGEMA_reg_buffer_11199 ( .C (clk), .D (new_AGEMA_signal_23922), .Q (new_AGEMA_signal_23923) ) ;
    buf_clk new_AGEMA_reg_buffer_11203 ( .C (clk), .D (new_AGEMA_signal_23926), .Q (new_AGEMA_signal_23927) ) ;
    buf_clk new_AGEMA_reg_buffer_11207 ( .C (clk), .D (new_AGEMA_signal_23930), .Q (new_AGEMA_signal_23931) ) ;
    buf_clk new_AGEMA_reg_buffer_11211 ( .C (clk), .D (new_AGEMA_signal_23934), .Q (new_AGEMA_signal_23935) ) ;
    buf_clk new_AGEMA_reg_buffer_11215 ( .C (clk), .D (new_AGEMA_signal_23938), .Q (new_AGEMA_signal_23939) ) ;
    buf_clk new_AGEMA_reg_buffer_11219 ( .C (clk), .D (new_AGEMA_signal_23942), .Q (new_AGEMA_signal_23943) ) ;
    buf_clk new_AGEMA_reg_buffer_11223 ( .C (clk), .D (new_AGEMA_signal_23946), .Q (new_AGEMA_signal_23947) ) ;
    buf_clk new_AGEMA_reg_buffer_11227 ( .C (clk), .D (new_AGEMA_signal_23950), .Q (new_AGEMA_signal_23951) ) ;
    buf_clk new_AGEMA_reg_buffer_11231 ( .C (clk), .D (new_AGEMA_signal_23954), .Q (new_AGEMA_signal_23955) ) ;
    buf_clk new_AGEMA_reg_buffer_11235 ( .C (clk), .D (new_AGEMA_signal_23958), .Q (new_AGEMA_signal_23959) ) ;
    buf_clk new_AGEMA_reg_buffer_11239 ( .C (clk), .D (new_AGEMA_signal_23962), .Q (new_AGEMA_signal_23963) ) ;
    buf_clk new_AGEMA_reg_buffer_11243 ( .C (clk), .D (new_AGEMA_signal_23966), .Q (new_AGEMA_signal_23967) ) ;
    buf_clk new_AGEMA_reg_buffer_11247 ( .C (clk), .D (new_AGEMA_signal_23970), .Q (new_AGEMA_signal_23971) ) ;
    buf_clk new_AGEMA_reg_buffer_11251 ( .C (clk), .D (new_AGEMA_signal_23974), .Q (new_AGEMA_signal_23975) ) ;
    buf_clk new_AGEMA_reg_buffer_11255 ( .C (clk), .D (new_AGEMA_signal_23978), .Q (new_AGEMA_signal_23979) ) ;
    buf_clk new_AGEMA_reg_buffer_11259 ( .C (clk), .D (new_AGEMA_signal_23982), .Q (new_AGEMA_signal_23983) ) ;
    buf_clk new_AGEMA_reg_buffer_11263 ( .C (clk), .D (new_AGEMA_signal_23986), .Q (new_AGEMA_signal_23987) ) ;
    buf_clk new_AGEMA_reg_buffer_11267 ( .C (clk), .D (new_AGEMA_signal_23990), .Q (new_AGEMA_signal_23991) ) ;
    buf_clk new_AGEMA_reg_buffer_11271 ( .C (clk), .D (new_AGEMA_signal_23994), .Q (new_AGEMA_signal_23995) ) ;
    buf_clk new_AGEMA_reg_buffer_11275 ( .C (clk), .D (new_AGEMA_signal_23998), .Q (new_AGEMA_signal_23999) ) ;
    buf_clk new_AGEMA_reg_buffer_11279 ( .C (clk), .D (new_AGEMA_signal_24002), .Q (new_AGEMA_signal_24003) ) ;
    buf_clk new_AGEMA_reg_buffer_11283 ( .C (clk), .D (new_AGEMA_signal_24006), .Q (new_AGEMA_signal_24007) ) ;
    buf_clk new_AGEMA_reg_buffer_11287 ( .C (clk), .D (new_AGEMA_signal_24010), .Q (new_AGEMA_signal_24011) ) ;
    buf_clk new_AGEMA_reg_buffer_11291 ( .C (clk), .D (new_AGEMA_signal_24014), .Q (new_AGEMA_signal_24015) ) ;
    buf_clk new_AGEMA_reg_buffer_11295 ( .C (clk), .D (new_AGEMA_signal_24018), .Q (new_AGEMA_signal_24019) ) ;
    buf_clk new_AGEMA_reg_buffer_11299 ( .C (clk), .D (new_AGEMA_signal_24022), .Q (new_AGEMA_signal_24023) ) ;
    buf_clk new_AGEMA_reg_buffer_11303 ( .C (clk), .D (new_AGEMA_signal_24026), .Q (new_AGEMA_signal_24027) ) ;
    buf_clk new_AGEMA_reg_buffer_11307 ( .C (clk), .D (new_AGEMA_signal_24030), .Q (new_AGEMA_signal_24031) ) ;
    buf_clk new_AGEMA_reg_buffer_11311 ( .C (clk), .D (new_AGEMA_signal_24034), .Q (new_AGEMA_signal_24035) ) ;
    buf_clk new_AGEMA_reg_buffer_11315 ( .C (clk), .D (new_AGEMA_signal_24038), .Q (new_AGEMA_signal_24039) ) ;
    buf_clk new_AGEMA_reg_buffer_11319 ( .C (clk), .D (new_AGEMA_signal_24042), .Q (new_AGEMA_signal_24043) ) ;
    buf_clk new_AGEMA_reg_buffer_11323 ( .C (clk), .D (new_AGEMA_signal_24046), .Q (new_AGEMA_signal_24047) ) ;
    buf_clk new_AGEMA_reg_buffer_11327 ( .C (clk), .D (new_AGEMA_signal_24050), .Q (new_AGEMA_signal_24051) ) ;
    buf_clk new_AGEMA_reg_buffer_11331 ( .C (clk), .D (new_AGEMA_signal_24054), .Q (new_AGEMA_signal_24055) ) ;
    buf_clk new_AGEMA_reg_buffer_11335 ( .C (clk), .D (new_AGEMA_signal_24058), .Q (new_AGEMA_signal_24059) ) ;
    buf_clk new_AGEMA_reg_buffer_11339 ( .C (clk), .D (new_AGEMA_signal_24062), .Q (new_AGEMA_signal_24063) ) ;
    buf_clk new_AGEMA_reg_buffer_11343 ( .C (clk), .D (new_AGEMA_signal_24066), .Q (new_AGEMA_signal_24067) ) ;
    buf_clk new_AGEMA_reg_buffer_11347 ( .C (clk), .D (new_AGEMA_signal_24070), .Q (new_AGEMA_signal_24071) ) ;
    buf_clk new_AGEMA_reg_buffer_11351 ( .C (clk), .D (new_AGEMA_signal_24074), .Q (new_AGEMA_signal_24075) ) ;
    buf_clk new_AGEMA_reg_buffer_11355 ( .C (clk), .D (new_AGEMA_signal_24078), .Q (new_AGEMA_signal_24079) ) ;
    buf_clk new_AGEMA_reg_buffer_11359 ( .C (clk), .D (new_AGEMA_signal_24082), .Q (new_AGEMA_signal_24083) ) ;
    buf_clk new_AGEMA_reg_buffer_11363 ( .C (clk), .D (new_AGEMA_signal_24086), .Q (new_AGEMA_signal_24087) ) ;
    buf_clk new_AGEMA_reg_buffer_11367 ( .C (clk), .D (new_AGEMA_signal_24090), .Q (new_AGEMA_signal_24091) ) ;
    buf_clk new_AGEMA_reg_buffer_11371 ( .C (clk), .D (new_AGEMA_signal_24094), .Q (new_AGEMA_signal_24095) ) ;
    buf_clk new_AGEMA_reg_buffer_11375 ( .C (clk), .D (new_AGEMA_signal_24098), .Q (new_AGEMA_signal_24099) ) ;
    buf_clk new_AGEMA_reg_buffer_11379 ( .C (clk), .D (new_AGEMA_signal_24102), .Q (new_AGEMA_signal_24103) ) ;
    buf_clk new_AGEMA_reg_buffer_11383 ( .C (clk), .D (new_AGEMA_signal_24106), .Q (new_AGEMA_signal_24107) ) ;
    buf_clk new_AGEMA_reg_buffer_11387 ( .C (clk), .D (new_AGEMA_signal_24110), .Q (new_AGEMA_signal_24111) ) ;
    buf_clk new_AGEMA_reg_buffer_11391 ( .C (clk), .D (new_AGEMA_signal_24114), .Q (new_AGEMA_signal_24115) ) ;
    buf_clk new_AGEMA_reg_buffer_11395 ( .C (clk), .D (new_AGEMA_signal_24118), .Q (new_AGEMA_signal_24119) ) ;
    buf_clk new_AGEMA_reg_buffer_11399 ( .C (clk), .D (new_AGEMA_signal_24122), .Q (new_AGEMA_signal_24123) ) ;
    buf_clk new_AGEMA_reg_buffer_11403 ( .C (clk), .D (new_AGEMA_signal_24126), .Q (new_AGEMA_signal_24127) ) ;
    buf_clk new_AGEMA_reg_buffer_11407 ( .C (clk), .D (new_AGEMA_signal_24130), .Q (new_AGEMA_signal_24131) ) ;
    buf_clk new_AGEMA_reg_buffer_11411 ( .C (clk), .D (new_AGEMA_signal_24134), .Q (new_AGEMA_signal_24135) ) ;
    buf_clk new_AGEMA_reg_buffer_11415 ( .C (clk), .D (new_AGEMA_signal_24138), .Q (new_AGEMA_signal_24139) ) ;
    buf_clk new_AGEMA_reg_buffer_11419 ( .C (clk), .D (new_AGEMA_signal_24142), .Q (new_AGEMA_signal_24143) ) ;
    buf_clk new_AGEMA_reg_buffer_11423 ( .C (clk), .D (new_AGEMA_signal_24146), .Q (new_AGEMA_signal_24147) ) ;
    buf_clk new_AGEMA_reg_buffer_11427 ( .C (clk), .D (new_AGEMA_signal_24150), .Q (new_AGEMA_signal_24151) ) ;
    buf_clk new_AGEMA_reg_buffer_11431 ( .C (clk), .D (new_AGEMA_signal_24154), .Q (new_AGEMA_signal_24155) ) ;
    buf_clk new_AGEMA_reg_buffer_11435 ( .C (clk), .D (new_AGEMA_signal_24158), .Q (new_AGEMA_signal_24159) ) ;
    buf_clk new_AGEMA_reg_buffer_11439 ( .C (clk), .D (new_AGEMA_signal_24162), .Q (new_AGEMA_signal_24163) ) ;
    buf_clk new_AGEMA_reg_buffer_11443 ( .C (clk), .D (new_AGEMA_signal_24166), .Q (new_AGEMA_signal_24167) ) ;
    buf_clk new_AGEMA_reg_buffer_11447 ( .C (clk), .D (new_AGEMA_signal_24170), .Q (new_AGEMA_signal_24171) ) ;
    buf_clk new_AGEMA_reg_buffer_11451 ( .C (clk), .D (new_AGEMA_signal_24174), .Q (new_AGEMA_signal_24175) ) ;
    buf_clk new_AGEMA_reg_buffer_11455 ( .C (clk), .D (new_AGEMA_signal_24178), .Q (new_AGEMA_signal_24179) ) ;
    buf_clk new_AGEMA_reg_buffer_11459 ( .C (clk), .D (new_AGEMA_signal_24182), .Q (new_AGEMA_signal_24183) ) ;
    buf_clk new_AGEMA_reg_buffer_11463 ( .C (clk), .D (new_AGEMA_signal_24186), .Q (new_AGEMA_signal_24187) ) ;
    buf_clk new_AGEMA_reg_buffer_11467 ( .C (clk), .D (new_AGEMA_signal_24190), .Q (new_AGEMA_signal_24191) ) ;
    buf_clk new_AGEMA_reg_buffer_11471 ( .C (clk), .D (new_AGEMA_signal_24194), .Q (new_AGEMA_signal_24195) ) ;
    buf_clk new_AGEMA_reg_buffer_11475 ( .C (clk), .D (new_AGEMA_signal_24198), .Q (new_AGEMA_signal_24199) ) ;
    buf_clk new_AGEMA_reg_buffer_11479 ( .C (clk), .D (new_AGEMA_signal_24202), .Q (new_AGEMA_signal_24203) ) ;
    buf_clk new_AGEMA_reg_buffer_11483 ( .C (clk), .D (new_AGEMA_signal_24206), .Q (new_AGEMA_signal_24207) ) ;
    buf_clk new_AGEMA_reg_buffer_11487 ( .C (clk), .D (new_AGEMA_signal_24210), .Q (new_AGEMA_signal_24211) ) ;
    buf_clk new_AGEMA_reg_buffer_11491 ( .C (clk), .D (new_AGEMA_signal_24214), .Q (new_AGEMA_signal_24215) ) ;
    buf_clk new_AGEMA_reg_buffer_11495 ( .C (clk), .D (new_AGEMA_signal_24218), .Q (new_AGEMA_signal_24219) ) ;
    buf_clk new_AGEMA_reg_buffer_11499 ( .C (clk), .D (new_AGEMA_signal_24222), .Q (new_AGEMA_signal_24223) ) ;
    buf_clk new_AGEMA_reg_buffer_11503 ( .C (clk), .D (new_AGEMA_signal_24226), .Q (new_AGEMA_signal_24227) ) ;
    buf_clk new_AGEMA_reg_buffer_11507 ( .C (clk), .D (new_AGEMA_signal_24230), .Q (new_AGEMA_signal_24231) ) ;
    buf_clk new_AGEMA_reg_buffer_11511 ( .C (clk), .D (new_AGEMA_signal_24234), .Q (new_AGEMA_signal_24235) ) ;
    buf_clk new_AGEMA_reg_buffer_11515 ( .C (clk), .D (new_AGEMA_signal_24238), .Q (new_AGEMA_signal_24239) ) ;
    buf_clk new_AGEMA_reg_buffer_11519 ( .C (clk), .D (new_AGEMA_signal_24242), .Q (new_AGEMA_signal_24243) ) ;
    buf_clk new_AGEMA_reg_buffer_11523 ( .C (clk), .D (new_AGEMA_signal_24246), .Q (new_AGEMA_signal_24247) ) ;
    buf_clk new_AGEMA_reg_buffer_11527 ( .C (clk), .D (new_AGEMA_signal_24250), .Q (new_AGEMA_signal_24251) ) ;
    buf_clk new_AGEMA_reg_buffer_11531 ( .C (clk), .D (new_AGEMA_signal_24254), .Q (new_AGEMA_signal_24255) ) ;
    buf_clk new_AGEMA_reg_buffer_11535 ( .C (clk), .D (new_AGEMA_signal_24258), .Q (new_AGEMA_signal_24259) ) ;
    buf_clk new_AGEMA_reg_buffer_11539 ( .C (clk), .D (new_AGEMA_signal_24262), .Q (new_AGEMA_signal_24263) ) ;
    buf_clk new_AGEMA_reg_buffer_11543 ( .C (clk), .D (new_AGEMA_signal_24266), .Q (new_AGEMA_signal_24267) ) ;
    buf_clk new_AGEMA_reg_buffer_11547 ( .C (clk), .D (new_AGEMA_signal_24270), .Q (new_AGEMA_signal_24271) ) ;
    buf_clk new_AGEMA_reg_buffer_11551 ( .C (clk), .D (new_AGEMA_signal_24274), .Q (new_AGEMA_signal_24275) ) ;
    buf_clk new_AGEMA_reg_buffer_11555 ( .C (clk), .D (new_AGEMA_signal_24278), .Q (new_AGEMA_signal_24279) ) ;
    buf_clk new_AGEMA_reg_buffer_11559 ( .C (clk), .D (new_AGEMA_signal_24282), .Q (new_AGEMA_signal_24283) ) ;
    buf_clk new_AGEMA_reg_buffer_11563 ( .C (clk), .D (new_AGEMA_signal_24286), .Q (new_AGEMA_signal_24287) ) ;
    buf_clk new_AGEMA_reg_buffer_11567 ( .C (clk), .D (new_AGEMA_signal_24290), .Q (new_AGEMA_signal_24291) ) ;
    buf_clk new_AGEMA_reg_buffer_11571 ( .C (clk), .D (new_AGEMA_signal_24294), .Q (new_AGEMA_signal_24295) ) ;
    buf_clk new_AGEMA_reg_buffer_11575 ( .C (clk), .D (new_AGEMA_signal_24298), .Q (new_AGEMA_signal_24299) ) ;
    buf_clk new_AGEMA_reg_buffer_11579 ( .C (clk), .D (new_AGEMA_signal_24302), .Q (new_AGEMA_signal_24303) ) ;
    buf_clk new_AGEMA_reg_buffer_11583 ( .C (clk), .D (new_AGEMA_signal_24306), .Q (new_AGEMA_signal_24307) ) ;
    buf_clk new_AGEMA_reg_buffer_11587 ( .C (clk), .D (new_AGEMA_signal_24310), .Q (new_AGEMA_signal_24311) ) ;
    buf_clk new_AGEMA_reg_buffer_11591 ( .C (clk), .D (new_AGEMA_signal_24314), .Q (new_AGEMA_signal_24315) ) ;
    buf_clk new_AGEMA_reg_buffer_11595 ( .C (clk), .D (new_AGEMA_signal_24318), .Q (new_AGEMA_signal_24319) ) ;
    buf_clk new_AGEMA_reg_buffer_11599 ( .C (clk), .D (new_AGEMA_signal_24322), .Q (new_AGEMA_signal_24323) ) ;
    buf_clk new_AGEMA_reg_buffer_11603 ( .C (clk), .D (new_AGEMA_signal_24326), .Q (new_AGEMA_signal_24327) ) ;
    buf_clk new_AGEMA_reg_buffer_11607 ( .C (clk), .D (new_AGEMA_signal_24330), .Q (new_AGEMA_signal_24331) ) ;
    buf_clk new_AGEMA_reg_buffer_11611 ( .C (clk), .D (new_AGEMA_signal_24334), .Q (new_AGEMA_signal_24335) ) ;
    buf_clk new_AGEMA_reg_buffer_11615 ( .C (clk), .D (new_AGEMA_signal_24338), .Q (new_AGEMA_signal_24339) ) ;
    buf_clk new_AGEMA_reg_buffer_11619 ( .C (clk), .D (new_AGEMA_signal_24342), .Q (new_AGEMA_signal_24343) ) ;
    buf_clk new_AGEMA_reg_buffer_11623 ( .C (clk), .D (new_AGEMA_signal_24346), .Q (new_AGEMA_signal_24347) ) ;
    buf_clk new_AGEMA_reg_buffer_11627 ( .C (clk), .D (new_AGEMA_signal_24350), .Q (new_AGEMA_signal_24351) ) ;
    buf_clk new_AGEMA_reg_buffer_11631 ( .C (clk), .D (new_AGEMA_signal_24354), .Q (new_AGEMA_signal_24355) ) ;
    buf_clk new_AGEMA_reg_buffer_11635 ( .C (clk), .D (new_AGEMA_signal_24358), .Q (new_AGEMA_signal_24359) ) ;
    buf_clk new_AGEMA_reg_buffer_11639 ( .C (clk), .D (new_AGEMA_signal_24362), .Q (new_AGEMA_signal_24363) ) ;
    buf_clk new_AGEMA_reg_buffer_11643 ( .C (clk), .D (new_AGEMA_signal_24366), .Q (new_AGEMA_signal_24367) ) ;
    buf_clk new_AGEMA_reg_buffer_11647 ( .C (clk), .D (new_AGEMA_signal_24370), .Q (new_AGEMA_signal_24371) ) ;
    buf_clk new_AGEMA_reg_buffer_11651 ( .C (clk), .D (new_AGEMA_signal_24374), .Q (new_AGEMA_signal_24375) ) ;
    buf_clk new_AGEMA_reg_buffer_11655 ( .C (clk), .D (new_AGEMA_signal_24378), .Q (new_AGEMA_signal_24379) ) ;
    buf_clk new_AGEMA_reg_buffer_11659 ( .C (clk), .D (new_AGEMA_signal_24382), .Q (new_AGEMA_signal_24383) ) ;
    buf_clk new_AGEMA_reg_buffer_11663 ( .C (clk), .D (new_AGEMA_signal_24386), .Q (new_AGEMA_signal_24387) ) ;
    buf_clk new_AGEMA_reg_buffer_11667 ( .C (clk), .D (new_AGEMA_signal_24390), .Q (new_AGEMA_signal_24391) ) ;
    buf_clk new_AGEMA_reg_buffer_11671 ( .C (clk), .D (new_AGEMA_signal_24394), .Q (new_AGEMA_signal_24395) ) ;
    buf_clk new_AGEMA_reg_buffer_11675 ( .C (clk), .D (new_AGEMA_signal_24398), .Q (new_AGEMA_signal_24399) ) ;
    buf_clk new_AGEMA_reg_buffer_11679 ( .C (clk), .D (new_AGEMA_signal_24402), .Q (new_AGEMA_signal_24403) ) ;
    buf_clk new_AGEMA_reg_buffer_11683 ( .C (clk), .D (new_AGEMA_signal_24406), .Q (new_AGEMA_signal_24407) ) ;
    buf_clk new_AGEMA_reg_buffer_11687 ( .C (clk), .D (new_AGEMA_signal_24410), .Q (new_AGEMA_signal_24411) ) ;
    buf_clk new_AGEMA_reg_buffer_11691 ( .C (clk), .D (new_AGEMA_signal_24414), .Q (new_AGEMA_signal_24415) ) ;
    buf_clk new_AGEMA_reg_buffer_11695 ( .C (clk), .D (new_AGEMA_signal_24418), .Q (new_AGEMA_signal_24419) ) ;
    buf_clk new_AGEMA_reg_buffer_11699 ( .C (clk), .D (new_AGEMA_signal_24422), .Q (new_AGEMA_signal_24423) ) ;
    buf_clk new_AGEMA_reg_buffer_11703 ( .C (clk), .D (new_AGEMA_signal_24426), .Q (new_AGEMA_signal_24427) ) ;
    buf_clk new_AGEMA_reg_buffer_11707 ( .C (clk), .D (new_AGEMA_signal_24430), .Q (new_AGEMA_signal_24431) ) ;
    buf_clk new_AGEMA_reg_buffer_11711 ( .C (clk), .D (new_AGEMA_signal_24434), .Q (new_AGEMA_signal_24435) ) ;
    buf_clk new_AGEMA_reg_buffer_11715 ( .C (clk), .D (new_AGEMA_signal_24438), .Q (new_AGEMA_signal_24439) ) ;
    buf_clk new_AGEMA_reg_buffer_11719 ( .C (clk), .D (new_AGEMA_signal_24442), .Q (new_AGEMA_signal_24443) ) ;
    buf_clk new_AGEMA_reg_buffer_11723 ( .C (clk), .D (new_AGEMA_signal_24446), .Q (new_AGEMA_signal_24447) ) ;
    buf_clk new_AGEMA_reg_buffer_11727 ( .C (clk), .D (new_AGEMA_signal_24450), .Q (new_AGEMA_signal_24451) ) ;
    buf_clk new_AGEMA_reg_buffer_11731 ( .C (clk), .D (new_AGEMA_signal_24454), .Q (new_AGEMA_signal_24455) ) ;
    buf_clk new_AGEMA_reg_buffer_11735 ( .C (clk), .D (new_AGEMA_signal_24458), .Q (new_AGEMA_signal_24459) ) ;
    buf_clk new_AGEMA_reg_buffer_11739 ( .C (clk), .D (new_AGEMA_signal_24462), .Q (new_AGEMA_signal_24463) ) ;
    buf_clk new_AGEMA_reg_buffer_11743 ( .C (clk), .D (new_AGEMA_signal_24466), .Q (new_AGEMA_signal_24467) ) ;
    buf_clk new_AGEMA_reg_buffer_11747 ( .C (clk), .D (new_AGEMA_signal_24470), .Q (new_AGEMA_signal_24471) ) ;
    buf_clk new_AGEMA_reg_buffer_11751 ( .C (clk), .D (new_AGEMA_signal_24474), .Q (new_AGEMA_signal_24475) ) ;
    buf_clk new_AGEMA_reg_buffer_11755 ( .C (clk), .D (new_AGEMA_signal_24478), .Q (new_AGEMA_signal_24479) ) ;
    buf_clk new_AGEMA_reg_buffer_11759 ( .C (clk), .D (new_AGEMA_signal_24482), .Q (new_AGEMA_signal_24483) ) ;
    buf_clk new_AGEMA_reg_buffer_11763 ( .C (clk), .D (new_AGEMA_signal_24486), .Q (new_AGEMA_signal_24487) ) ;
    buf_clk new_AGEMA_reg_buffer_11767 ( .C (clk), .D (new_AGEMA_signal_24490), .Q (new_AGEMA_signal_24491) ) ;
    buf_clk new_AGEMA_reg_buffer_11771 ( .C (clk), .D (new_AGEMA_signal_24494), .Q (new_AGEMA_signal_24495) ) ;
    buf_clk new_AGEMA_reg_buffer_11775 ( .C (clk), .D (new_AGEMA_signal_24498), .Q (new_AGEMA_signal_24499) ) ;
    buf_clk new_AGEMA_reg_buffer_11779 ( .C (clk), .D (new_AGEMA_signal_24502), .Q (new_AGEMA_signal_24503) ) ;
    buf_clk new_AGEMA_reg_buffer_11783 ( .C (clk), .D (new_AGEMA_signal_24506), .Q (new_AGEMA_signal_24507) ) ;
    buf_clk new_AGEMA_reg_buffer_11787 ( .C (clk), .D (new_AGEMA_signal_24510), .Q (new_AGEMA_signal_24511) ) ;
    buf_clk new_AGEMA_reg_buffer_11791 ( .C (clk), .D (new_AGEMA_signal_24514), .Q (new_AGEMA_signal_24515) ) ;
    buf_clk new_AGEMA_reg_buffer_11795 ( .C (clk), .D (new_AGEMA_signal_24518), .Q (new_AGEMA_signal_24519) ) ;
    buf_clk new_AGEMA_reg_buffer_11799 ( .C (clk), .D (new_AGEMA_signal_24522), .Q (new_AGEMA_signal_24523) ) ;
    buf_clk new_AGEMA_reg_buffer_11803 ( .C (clk), .D (new_AGEMA_signal_24526), .Q (new_AGEMA_signal_24527) ) ;
    buf_clk new_AGEMA_reg_buffer_11807 ( .C (clk), .D (new_AGEMA_signal_24530), .Q (new_AGEMA_signal_24531) ) ;
    buf_clk new_AGEMA_reg_buffer_11811 ( .C (clk), .D (new_AGEMA_signal_24534), .Q (new_AGEMA_signal_24535) ) ;
    buf_clk new_AGEMA_reg_buffer_11815 ( .C (clk), .D (new_AGEMA_signal_24538), .Q (new_AGEMA_signal_24539) ) ;
    buf_clk new_AGEMA_reg_buffer_11819 ( .C (clk), .D (new_AGEMA_signal_24542), .Q (new_AGEMA_signal_24543) ) ;
    buf_clk new_AGEMA_reg_buffer_11823 ( .C (clk), .D (new_AGEMA_signal_24546), .Q (new_AGEMA_signal_24547) ) ;
    buf_clk new_AGEMA_reg_buffer_11827 ( .C (clk), .D (new_AGEMA_signal_24550), .Q (new_AGEMA_signal_24551) ) ;
    buf_clk new_AGEMA_reg_buffer_11831 ( .C (clk), .D (new_AGEMA_signal_24554), .Q (new_AGEMA_signal_24555) ) ;
    buf_clk new_AGEMA_reg_buffer_11835 ( .C (clk), .D (new_AGEMA_signal_24558), .Q (new_AGEMA_signal_24559) ) ;
    buf_clk new_AGEMA_reg_buffer_11839 ( .C (clk), .D (new_AGEMA_signal_24562), .Q (new_AGEMA_signal_24563) ) ;
    buf_clk new_AGEMA_reg_buffer_11843 ( .C (clk), .D (new_AGEMA_signal_24566), .Q (new_AGEMA_signal_24567) ) ;
    buf_clk new_AGEMA_reg_buffer_11847 ( .C (clk), .D (new_AGEMA_signal_24570), .Q (new_AGEMA_signal_24571) ) ;
    buf_clk new_AGEMA_reg_buffer_11851 ( .C (clk), .D (new_AGEMA_signal_24574), .Q (new_AGEMA_signal_24575) ) ;
    buf_clk new_AGEMA_reg_buffer_11855 ( .C (clk), .D (new_AGEMA_signal_24578), .Q (new_AGEMA_signal_24579) ) ;
    buf_clk new_AGEMA_reg_buffer_11859 ( .C (clk), .D (new_AGEMA_signal_24582), .Q (new_AGEMA_signal_24583) ) ;
    buf_clk new_AGEMA_reg_buffer_11863 ( .C (clk), .D (new_AGEMA_signal_24586), .Q (new_AGEMA_signal_24587) ) ;
    buf_clk new_AGEMA_reg_buffer_11867 ( .C (clk), .D (new_AGEMA_signal_24590), .Q (new_AGEMA_signal_24591) ) ;
    buf_clk new_AGEMA_reg_buffer_11871 ( .C (clk), .D (new_AGEMA_signal_24594), .Q (new_AGEMA_signal_24595) ) ;
    buf_clk new_AGEMA_reg_buffer_11875 ( .C (clk), .D (new_AGEMA_signal_24598), .Q (new_AGEMA_signal_24599) ) ;
    buf_clk new_AGEMA_reg_buffer_11879 ( .C (clk), .D (new_AGEMA_signal_24602), .Q (new_AGEMA_signal_24603) ) ;
    buf_clk new_AGEMA_reg_buffer_11883 ( .C (clk), .D (new_AGEMA_signal_24606), .Q (new_AGEMA_signal_24607) ) ;
    buf_clk new_AGEMA_reg_buffer_11887 ( .C (clk), .D (new_AGEMA_signal_24610), .Q (new_AGEMA_signal_24611) ) ;
    buf_clk new_AGEMA_reg_buffer_11891 ( .C (clk), .D (new_AGEMA_signal_24614), .Q (new_AGEMA_signal_24615) ) ;
    buf_clk new_AGEMA_reg_buffer_11895 ( .C (clk), .D (new_AGEMA_signal_24618), .Q (new_AGEMA_signal_24619) ) ;
    buf_clk new_AGEMA_reg_buffer_11899 ( .C (clk), .D (new_AGEMA_signal_24622), .Q (new_AGEMA_signal_24623) ) ;
    buf_clk new_AGEMA_reg_buffer_11903 ( .C (clk), .D (new_AGEMA_signal_24626), .Q (new_AGEMA_signal_24627) ) ;
    buf_clk new_AGEMA_reg_buffer_11907 ( .C (clk), .D (new_AGEMA_signal_24630), .Q (new_AGEMA_signal_24631) ) ;
    buf_clk new_AGEMA_reg_buffer_11911 ( .C (clk), .D (new_AGEMA_signal_24634), .Q (new_AGEMA_signal_24635) ) ;
    buf_clk new_AGEMA_reg_buffer_11915 ( .C (clk), .D (new_AGEMA_signal_24638), .Q (new_AGEMA_signal_24639) ) ;
    buf_clk new_AGEMA_reg_buffer_11919 ( .C (clk), .D (new_AGEMA_signal_24642), .Q (new_AGEMA_signal_24643) ) ;
    buf_clk new_AGEMA_reg_buffer_11923 ( .C (clk), .D (new_AGEMA_signal_24646), .Q (new_AGEMA_signal_24647) ) ;
    buf_clk new_AGEMA_reg_buffer_11927 ( .C (clk), .D (new_AGEMA_signal_24650), .Q (new_AGEMA_signal_24651) ) ;
    buf_clk new_AGEMA_reg_buffer_11931 ( .C (clk), .D (new_AGEMA_signal_24654), .Q (new_AGEMA_signal_24655) ) ;
    buf_clk new_AGEMA_reg_buffer_11935 ( .C (clk), .D (new_AGEMA_signal_24658), .Q (new_AGEMA_signal_24659) ) ;
    buf_clk new_AGEMA_reg_buffer_11939 ( .C (clk), .D (new_AGEMA_signal_24662), .Q (new_AGEMA_signal_24663) ) ;
    buf_clk new_AGEMA_reg_buffer_11943 ( .C (clk), .D (new_AGEMA_signal_24666), .Q (new_AGEMA_signal_24667) ) ;
    buf_clk new_AGEMA_reg_buffer_11947 ( .C (clk), .D (new_AGEMA_signal_24670), .Q (new_AGEMA_signal_24671) ) ;
    buf_clk new_AGEMA_reg_buffer_11951 ( .C (clk), .D (new_AGEMA_signal_24674), .Q (new_AGEMA_signal_24675) ) ;
    buf_clk new_AGEMA_reg_buffer_11955 ( .C (clk), .D (new_AGEMA_signal_24678), .Q (new_AGEMA_signal_24679) ) ;
    buf_clk new_AGEMA_reg_buffer_11959 ( .C (clk), .D (new_AGEMA_signal_24682), .Q (new_AGEMA_signal_24683) ) ;
    buf_clk new_AGEMA_reg_buffer_11963 ( .C (clk), .D (new_AGEMA_signal_24686), .Q (new_AGEMA_signal_24687) ) ;
    buf_clk new_AGEMA_reg_buffer_11967 ( .C (clk), .D (new_AGEMA_signal_24690), .Q (new_AGEMA_signal_24691) ) ;
    buf_clk new_AGEMA_reg_buffer_11971 ( .C (clk), .D (new_AGEMA_signal_24694), .Q (new_AGEMA_signal_24695) ) ;
    buf_clk new_AGEMA_reg_buffer_11975 ( .C (clk), .D (new_AGEMA_signal_24698), .Q (new_AGEMA_signal_24699) ) ;
    buf_clk new_AGEMA_reg_buffer_11979 ( .C (clk), .D (new_AGEMA_signal_24702), .Q (new_AGEMA_signal_24703) ) ;
    buf_clk new_AGEMA_reg_buffer_11983 ( .C (clk), .D (new_AGEMA_signal_24706), .Q (new_AGEMA_signal_24707) ) ;
    buf_clk new_AGEMA_reg_buffer_11987 ( .C (clk), .D (new_AGEMA_signal_24710), .Q (new_AGEMA_signal_24711) ) ;
    buf_clk new_AGEMA_reg_buffer_11991 ( .C (clk), .D (new_AGEMA_signal_24714), .Q (new_AGEMA_signal_24715) ) ;
    buf_clk new_AGEMA_reg_buffer_11995 ( .C (clk), .D (new_AGEMA_signal_24718), .Q (new_AGEMA_signal_24719) ) ;
    buf_clk new_AGEMA_reg_buffer_11999 ( .C (clk), .D (new_AGEMA_signal_24722), .Q (new_AGEMA_signal_24723) ) ;
    buf_clk new_AGEMA_reg_buffer_12003 ( .C (clk), .D (new_AGEMA_signal_24726), .Q (new_AGEMA_signal_24727) ) ;
    buf_clk new_AGEMA_reg_buffer_12007 ( .C (clk), .D (new_AGEMA_signal_24730), .Q (new_AGEMA_signal_24731) ) ;
    buf_clk new_AGEMA_reg_buffer_12011 ( .C (clk), .D (new_AGEMA_signal_24734), .Q (new_AGEMA_signal_24735) ) ;
    buf_clk new_AGEMA_reg_buffer_12015 ( .C (clk), .D (new_AGEMA_signal_24738), .Q (new_AGEMA_signal_24739) ) ;
    buf_clk new_AGEMA_reg_buffer_12019 ( .C (clk), .D (new_AGEMA_signal_24742), .Q (new_AGEMA_signal_24743) ) ;
    buf_clk new_AGEMA_reg_buffer_12023 ( .C (clk), .D (new_AGEMA_signal_24746), .Q (new_AGEMA_signal_24747) ) ;
    buf_clk new_AGEMA_reg_buffer_12027 ( .C (clk), .D (new_AGEMA_signal_24750), .Q (new_AGEMA_signal_24751) ) ;
    buf_clk new_AGEMA_reg_buffer_12031 ( .C (clk), .D (new_AGEMA_signal_24754), .Q (new_AGEMA_signal_24755) ) ;
    buf_clk new_AGEMA_reg_buffer_12035 ( .C (clk), .D (new_AGEMA_signal_24758), .Q (new_AGEMA_signal_24759) ) ;
    buf_clk new_AGEMA_reg_buffer_12039 ( .C (clk), .D (new_AGEMA_signal_24762), .Q (new_AGEMA_signal_24763) ) ;
    buf_clk new_AGEMA_reg_buffer_12043 ( .C (clk), .D (new_AGEMA_signal_24766), .Q (new_AGEMA_signal_24767) ) ;
    buf_clk new_AGEMA_reg_buffer_12047 ( .C (clk), .D (new_AGEMA_signal_24770), .Q (new_AGEMA_signal_24771) ) ;
    buf_clk new_AGEMA_reg_buffer_12051 ( .C (clk), .D (new_AGEMA_signal_24774), .Q (new_AGEMA_signal_24775) ) ;
    buf_clk new_AGEMA_reg_buffer_12055 ( .C (clk), .D (new_AGEMA_signal_24778), .Q (new_AGEMA_signal_24779) ) ;
    buf_clk new_AGEMA_reg_buffer_12059 ( .C (clk), .D (new_AGEMA_signal_24782), .Q (new_AGEMA_signal_24783) ) ;
    buf_clk new_AGEMA_reg_buffer_12063 ( .C (clk), .D (new_AGEMA_signal_24786), .Q (new_AGEMA_signal_24787) ) ;
    buf_clk new_AGEMA_reg_buffer_12067 ( .C (clk), .D (new_AGEMA_signal_24790), .Q (new_AGEMA_signal_24791) ) ;
    buf_clk new_AGEMA_reg_buffer_12071 ( .C (clk), .D (new_AGEMA_signal_24794), .Q (new_AGEMA_signal_24795) ) ;
    buf_clk new_AGEMA_reg_buffer_12075 ( .C (clk), .D (new_AGEMA_signal_24798), .Q (new_AGEMA_signal_24799) ) ;
    buf_clk new_AGEMA_reg_buffer_12079 ( .C (clk), .D (new_AGEMA_signal_24802), .Q (new_AGEMA_signal_24803) ) ;
    buf_clk new_AGEMA_reg_buffer_12083 ( .C (clk), .D (new_AGEMA_signal_24806), .Q (new_AGEMA_signal_24807) ) ;
    buf_clk new_AGEMA_reg_buffer_12087 ( .C (clk), .D (new_AGEMA_signal_24810), .Q (new_AGEMA_signal_24811) ) ;
    buf_clk new_AGEMA_reg_buffer_12091 ( .C (clk), .D (new_AGEMA_signal_24814), .Q (new_AGEMA_signal_24815) ) ;
    buf_clk new_AGEMA_reg_buffer_12095 ( .C (clk), .D (new_AGEMA_signal_24818), .Q (new_AGEMA_signal_24819) ) ;
    buf_clk new_AGEMA_reg_buffer_12099 ( .C (clk), .D (new_AGEMA_signal_24822), .Q (new_AGEMA_signal_24823) ) ;
    buf_clk new_AGEMA_reg_buffer_12103 ( .C (clk), .D (new_AGEMA_signal_24826), .Q (new_AGEMA_signal_24827) ) ;
    buf_clk new_AGEMA_reg_buffer_12107 ( .C (clk), .D (new_AGEMA_signal_24830), .Q (new_AGEMA_signal_24831) ) ;
    buf_clk new_AGEMA_reg_buffer_12111 ( .C (clk), .D (new_AGEMA_signal_24834), .Q (new_AGEMA_signal_24835) ) ;
    buf_clk new_AGEMA_reg_buffer_12115 ( .C (clk), .D (new_AGEMA_signal_24838), .Q (new_AGEMA_signal_24839) ) ;
    buf_clk new_AGEMA_reg_buffer_12119 ( .C (clk), .D (new_AGEMA_signal_24842), .Q (new_AGEMA_signal_24843) ) ;
    buf_clk new_AGEMA_reg_buffer_12123 ( .C (clk), .D (new_AGEMA_signal_24846), .Q (new_AGEMA_signal_24847) ) ;
    buf_clk new_AGEMA_reg_buffer_12127 ( .C (clk), .D (new_AGEMA_signal_24850), .Q (new_AGEMA_signal_24851) ) ;
    buf_clk new_AGEMA_reg_buffer_12131 ( .C (clk), .D (new_AGEMA_signal_24854), .Q (new_AGEMA_signal_24855) ) ;
    buf_clk new_AGEMA_reg_buffer_12135 ( .C (clk), .D (new_AGEMA_signal_24858), .Q (new_AGEMA_signal_24859) ) ;
    buf_clk new_AGEMA_reg_buffer_12139 ( .C (clk), .D (new_AGEMA_signal_24862), .Q (new_AGEMA_signal_24863) ) ;
    buf_clk new_AGEMA_reg_buffer_12143 ( .C (clk), .D (new_AGEMA_signal_24866), .Q (new_AGEMA_signal_24867) ) ;
    buf_clk new_AGEMA_reg_buffer_12147 ( .C (clk), .D (new_AGEMA_signal_24870), .Q (new_AGEMA_signal_24871) ) ;
    buf_clk new_AGEMA_reg_buffer_12151 ( .C (clk), .D (new_AGEMA_signal_24874), .Q (new_AGEMA_signal_24875) ) ;
    buf_clk new_AGEMA_reg_buffer_12155 ( .C (clk), .D (new_AGEMA_signal_24878), .Q (new_AGEMA_signal_24879) ) ;
    buf_clk new_AGEMA_reg_buffer_12159 ( .C (clk), .D (new_AGEMA_signal_24882), .Q (new_AGEMA_signal_24883) ) ;
    buf_clk new_AGEMA_reg_buffer_12163 ( .C (clk), .D (new_AGEMA_signal_24886), .Q (new_AGEMA_signal_24887) ) ;
    buf_clk new_AGEMA_reg_buffer_12167 ( .C (clk), .D (new_AGEMA_signal_24890), .Q (new_AGEMA_signal_24891) ) ;
    buf_clk new_AGEMA_reg_buffer_12171 ( .C (clk), .D (new_AGEMA_signal_24894), .Q (new_AGEMA_signal_24895) ) ;
    buf_clk new_AGEMA_reg_buffer_12175 ( .C (clk), .D (new_AGEMA_signal_24898), .Q (new_AGEMA_signal_24899) ) ;
    buf_clk new_AGEMA_reg_buffer_12179 ( .C (clk), .D (new_AGEMA_signal_24902), .Q (new_AGEMA_signal_24903) ) ;
    buf_clk new_AGEMA_reg_buffer_12183 ( .C (clk), .D (new_AGEMA_signal_24906), .Q (new_AGEMA_signal_24907) ) ;
    buf_clk new_AGEMA_reg_buffer_12187 ( .C (clk), .D (new_AGEMA_signal_24910), .Q (new_AGEMA_signal_24911) ) ;
    buf_clk new_AGEMA_reg_buffer_12191 ( .C (clk), .D (new_AGEMA_signal_24914), .Q (new_AGEMA_signal_24915) ) ;
    buf_clk new_AGEMA_reg_buffer_12195 ( .C (clk), .D (new_AGEMA_signal_24918), .Q (new_AGEMA_signal_24919) ) ;
    buf_clk new_AGEMA_reg_buffer_12198 ( .C (clk), .D (new_AGEMA_signal_24921), .Q (new_AGEMA_signal_24922) ) ;
    buf_clk new_AGEMA_reg_buffer_12201 ( .C (clk), .D (new_AGEMA_signal_24924), .Q (new_AGEMA_signal_24925) ) ;
    buf_clk new_AGEMA_reg_buffer_12204 ( .C (clk), .D (new_AGEMA_signal_24927), .Q (new_AGEMA_signal_24928) ) ;
    buf_clk new_AGEMA_reg_buffer_12207 ( .C (clk), .D (new_AGEMA_signal_24930), .Q (new_AGEMA_signal_24931) ) ;
    buf_clk new_AGEMA_reg_buffer_12210 ( .C (clk), .D (new_AGEMA_signal_24933), .Q (new_AGEMA_signal_24934) ) ;
    buf_clk new_AGEMA_reg_buffer_12213 ( .C (clk), .D (new_AGEMA_signal_24936), .Q (new_AGEMA_signal_24937) ) ;
    buf_clk new_AGEMA_reg_buffer_12216 ( .C (clk), .D (new_AGEMA_signal_24939), .Q (new_AGEMA_signal_24940) ) ;
    buf_clk new_AGEMA_reg_buffer_12219 ( .C (clk), .D (new_AGEMA_signal_24942), .Q (new_AGEMA_signal_24943) ) ;
    buf_clk new_AGEMA_reg_buffer_12222 ( .C (clk), .D (new_AGEMA_signal_24945), .Q (new_AGEMA_signal_24946) ) ;
    buf_clk new_AGEMA_reg_buffer_12225 ( .C (clk), .D (new_AGEMA_signal_24948), .Q (new_AGEMA_signal_24949) ) ;
    buf_clk new_AGEMA_reg_buffer_12228 ( .C (clk), .D (new_AGEMA_signal_24951), .Q (new_AGEMA_signal_24952) ) ;
    buf_clk new_AGEMA_reg_buffer_12231 ( .C (clk), .D (new_AGEMA_signal_24954), .Q (new_AGEMA_signal_24955) ) ;
    buf_clk new_AGEMA_reg_buffer_12234 ( .C (clk), .D (new_AGEMA_signal_24957), .Q (new_AGEMA_signal_24958) ) ;
    buf_clk new_AGEMA_reg_buffer_12237 ( .C (clk), .D (new_AGEMA_signal_24960), .Q (new_AGEMA_signal_24961) ) ;
    buf_clk new_AGEMA_reg_buffer_12240 ( .C (clk), .D (new_AGEMA_signal_24963), .Q (new_AGEMA_signal_24964) ) ;
    buf_clk new_AGEMA_reg_buffer_12243 ( .C (clk), .D (new_AGEMA_signal_24966), .Q (new_AGEMA_signal_24967) ) ;
    buf_clk new_AGEMA_reg_buffer_12246 ( .C (clk), .D (new_AGEMA_signal_24969), .Q (new_AGEMA_signal_24970) ) ;
    buf_clk new_AGEMA_reg_buffer_12249 ( .C (clk), .D (new_AGEMA_signal_24972), .Q (new_AGEMA_signal_24973) ) ;
    buf_clk new_AGEMA_reg_buffer_12252 ( .C (clk), .D (new_AGEMA_signal_24975), .Q (new_AGEMA_signal_24976) ) ;
    buf_clk new_AGEMA_reg_buffer_12255 ( .C (clk), .D (new_AGEMA_signal_24978), .Q (new_AGEMA_signal_24979) ) ;
    buf_clk new_AGEMA_reg_buffer_12258 ( .C (clk), .D (new_AGEMA_signal_24981), .Q (new_AGEMA_signal_24982) ) ;
    buf_clk new_AGEMA_reg_buffer_12261 ( .C (clk), .D (new_AGEMA_signal_24984), .Q (new_AGEMA_signal_24985) ) ;
    buf_clk new_AGEMA_reg_buffer_12264 ( .C (clk), .D (new_AGEMA_signal_24987), .Q (new_AGEMA_signal_24988) ) ;
    buf_clk new_AGEMA_reg_buffer_12267 ( .C (clk), .D (new_AGEMA_signal_24990), .Q (new_AGEMA_signal_24991) ) ;
    buf_clk new_AGEMA_reg_buffer_12270 ( .C (clk), .D (new_AGEMA_signal_24993), .Q (new_AGEMA_signal_24994) ) ;
    buf_clk new_AGEMA_reg_buffer_12273 ( .C (clk), .D (new_AGEMA_signal_24996), .Q (new_AGEMA_signal_24997) ) ;
    buf_clk new_AGEMA_reg_buffer_12276 ( .C (clk), .D (new_AGEMA_signal_24999), .Q (new_AGEMA_signal_25000) ) ;
    buf_clk new_AGEMA_reg_buffer_12279 ( .C (clk), .D (new_AGEMA_signal_25002), .Q (new_AGEMA_signal_25003) ) ;
    buf_clk new_AGEMA_reg_buffer_12282 ( .C (clk), .D (new_AGEMA_signal_25005), .Q (new_AGEMA_signal_25006) ) ;
    buf_clk new_AGEMA_reg_buffer_12285 ( .C (clk), .D (new_AGEMA_signal_25008), .Q (new_AGEMA_signal_25009) ) ;
    buf_clk new_AGEMA_reg_buffer_12288 ( .C (clk), .D (new_AGEMA_signal_25011), .Q (new_AGEMA_signal_25012) ) ;
    buf_clk new_AGEMA_reg_buffer_12291 ( .C (clk), .D (new_AGEMA_signal_25014), .Q (new_AGEMA_signal_25015) ) ;
    buf_clk new_AGEMA_reg_buffer_12294 ( .C (clk), .D (new_AGEMA_signal_25017), .Q (new_AGEMA_signal_25018) ) ;
    buf_clk new_AGEMA_reg_buffer_12297 ( .C (clk), .D (new_AGEMA_signal_25020), .Q (new_AGEMA_signal_25021) ) ;
    buf_clk new_AGEMA_reg_buffer_12300 ( .C (clk), .D (new_AGEMA_signal_25023), .Q (new_AGEMA_signal_25024) ) ;
    buf_clk new_AGEMA_reg_buffer_12303 ( .C (clk), .D (new_AGEMA_signal_25026), .Q (new_AGEMA_signal_25027) ) ;
    buf_clk new_AGEMA_reg_buffer_12306 ( .C (clk), .D (new_AGEMA_signal_25029), .Q (new_AGEMA_signal_25030) ) ;
    buf_clk new_AGEMA_reg_buffer_12309 ( .C (clk), .D (new_AGEMA_signal_25032), .Q (new_AGEMA_signal_25033) ) ;
    buf_clk new_AGEMA_reg_buffer_12312 ( .C (clk), .D (new_AGEMA_signal_25035), .Q (new_AGEMA_signal_25036) ) ;
    buf_clk new_AGEMA_reg_buffer_12315 ( .C (clk), .D (new_AGEMA_signal_25038), .Q (new_AGEMA_signal_25039) ) ;
    buf_clk new_AGEMA_reg_buffer_12318 ( .C (clk), .D (new_AGEMA_signal_25041), .Q (new_AGEMA_signal_25042) ) ;
    buf_clk new_AGEMA_reg_buffer_12321 ( .C (clk), .D (new_AGEMA_signal_25044), .Q (new_AGEMA_signal_25045) ) ;
    buf_clk new_AGEMA_reg_buffer_12324 ( .C (clk), .D (new_AGEMA_signal_25047), .Q (new_AGEMA_signal_25048) ) ;
    buf_clk new_AGEMA_reg_buffer_12327 ( .C (clk), .D (new_AGEMA_signal_25050), .Q (new_AGEMA_signal_25051) ) ;
    buf_clk new_AGEMA_reg_buffer_12330 ( .C (clk), .D (new_AGEMA_signal_25053), .Q (new_AGEMA_signal_25054) ) ;
    buf_clk new_AGEMA_reg_buffer_12333 ( .C (clk), .D (new_AGEMA_signal_25056), .Q (new_AGEMA_signal_25057) ) ;
    buf_clk new_AGEMA_reg_buffer_12336 ( .C (clk), .D (new_AGEMA_signal_25059), .Q (new_AGEMA_signal_25060) ) ;
    buf_clk new_AGEMA_reg_buffer_12339 ( .C (clk), .D (new_AGEMA_signal_25062), .Q (new_AGEMA_signal_25063) ) ;
    buf_clk new_AGEMA_reg_buffer_12342 ( .C (clk), .D (new_AGEMA_signal_25065), .Q (new_AGEMA_signal_25066) ) ;
    buf_clk new_AGEMA_reg_buffer_12345 ( .C (clk), .D (new_AGEMA_signal_25068), .Q (new_AGEMA_signal_25069) ) ;
    buf_clk new_AGEMA_reg_buffer_12348 ( .C (clk), .D (new_AGEMA_signal_25071), .Q (new_AGEMA_signal_25072) ) ;
    buf_clk new_AGEMA_reg_buffer_12351 ( .C (clk), .D (new_AGEMA_signal_25074), .Q (new_AGEMA_signal_25075) ) ;
    buf_clk new_AGEMA_reg_buffer_12354 ( .C (clk), .D (new_AGEMA_signal_25077), .Q (new_AGEMA_signal_25078) ) ;
    buf_clk new_AGEMA_reg_buffer_12357 ( .C (clk), .D (new_AGEMA_signal_25080), .Q (new_AGEMA_signal_25081) ) ;
    buf_clk new_AGEMA_reg_buffer_12360 ( .C (clk), .D (new_AGEMA_signal_25083), .Q (new_AGEMA_signal_25084) ) ;
    buf_clk new_AGEMA_reg_buffer_12363 ( .C (clk), .D (new_AGEMA_signal_25086), .Q (new_AGEMA_signal_25087) ) ;
    buf_clk new_AGEMA_reg_buffer_12366 ( .C (clk), .D (new_AGEMA_signal_25089), .Q (new_AGEMA_signal_25090) ) ;
    buf_clk new_AGEMA_reg_buffer_12369 ( .C (clk), .D (new_AGEMA_signal_25092), .Q (new_AGEMA_signal_25093) ) ;
    buf_clk new_AGEMA_reg_buffer_12372 ( .C (clk), .D (new_AGEMA_signal_25095), .Q (new_AGEMA_signal_25096) ) ;
    buf_clk new_AGEMA_reg_buffer_12375 ( .C (clk), .D (new_AGEMA_signal_25098), .Q (new_AGEMA_signal_25099) ) ;
    buf_clk new_AGEMA_reg_buffer_12378 ( .C (clk), .D (new_AGEMA_signal_25101), .Q (new_AGEMA_signal_25102) ) ;
    buf_clk new_AGEMA_reg_buffer_12381 ( .C (clk), .D (new_AGEMA_signal_25104), .Q (new_AGEMA_signal_25105) ) ;
    buf_clk new_AGEMA_reg_buffer_12384 ( .C (clk), .D (new_AGEMA_signal_25107), .Q (new_AGEMA_signal_25108) ) ;
    buf_clk new_AGEMA_reg_buffer_12387 ( .C (clk), .D (new_AGEMA_signal_25110), .Q (new_AGEMA_signal_25111) ) ;
    buf_clk new_AGEMA_reg_buffer_12390 ( .C (clk), .D (new_AGEMA_signal_25113), .Q (new_AGEMA_signal_25114) ) ;
    buf_clk new_AGEMA_reg_buffer_12393 ( .C (clk), .D (new_AGEMA_signal_25116), .Q (new_AGEMA_signal_25117) ) ;
    buf_clk new_AGEMA_reg_buffer_12396 ( .C (clk), .D (new_AGEMA_signal_25119), .Q (new_AGEMA_signal_25120) ) ;
    buf_clk new_AGEMA_reg_buffer_12399 ( .C (clk), .D (new_AGEMA_signal_25122), .Q (new_AGEMA_signal_25123) ) ;
    buf_clk new_AGEMA_reg_buffer_12402 ( .C (clk), .D (new_AGEMA_signal_25125), .Q (new_AGEMA_signal_25126) ) ;
    buf_clk new_AGEMA_reg_buffer_12405 ( .C (clk), .D (new_AGEMA_signal_25128), .Q (new_AGEMA_signal_25129) ) ;
    buf_clk new_AGEMA_reg_buffer_12408 ( .C (clk), .D (new_AGEMA_signal_25131), .Q (new_AGEMA_signal_25132) ) ;
    buf_clk new_AGEMA_reg_buffer_12411 ( .C (clk), .D (new_AGEMA_signal_25134), .Q (new_AGEMA_signal_25135) ) ;
    buf_clk new_AGEMA_reg_buffer_12414 ( .C (clk), .D (new_AGEMA_signal_25137), .Q (new_AGEMA_signal_25138) ) ;
    buf_clk new_AGEMA_reg_buffer_12417 ( .C (clk), .D (new_AGEMA_signal_25140), .Q (new_AGEMA_signal_25141) ) ;
    buf_clk new_AGEMA_reg_buffer_12420 ( .C (clk), .D (new_AGEMA_signal_25143), .Q (new_AGEMA_signal_25144) ) ;
    buf_clk new_AGEMA_reg_buffer_12423 ( .C (clk), .D (new_AGEMA_signal_25146), .Q (new_AGEMA_signal_25147) ) ;
    buf_clk new_AGEMA_reg_buffer_12426 ( .C (clk), .D (new_AGEMA_signal_25149), .Q (new_AGEMA_signal_25150) ) ;
    buf_clk new_AGEMA_reg_buffer_12429 ( .C (clk), .D (new_AGEMA_signal_25152), .Q (new_AGEMA_signal_25153) ) ;
    buf_clk new_AGEMA_reg_buffer_12432 ( .C (clk), .D (new_AGEMA_signal_25155), .Q (new_AGEMA_signal_25156) ) ;
    buf_clk new_AGEMA_reg_buffer_12435 ( .C (clk), .D (new_AGEMA_signal_25158), .Q (new_AGEMA_signal_25159) ) ;
    buf_clk new_AGEMA_reg_buffer_12438 ( .C (clk), .D (new_AGEMA_signal_25161), .Q (new_AGEMA_signal_25162) ) ;
    buf_clk new_AGEMA_reg_buffer_12441 ( .C (clk), .D (new_AGEMA_signal_25164), .Q (new_AGEMA_signal_25165) ) ;
    buf_clk new_AGEMA_reg_buffer_12444 ( .C (clk), .D (new_AGEMA_signal_25167), .Q (new_AGEMA_signal_25168) ) ;
    buf_clk new_AGEMA_reg_buffer_12447 ( .C (clk), .D (new_AGEMA_signal_25170), .Q (new_AGEMA_signal_25171) ) ;
    buf_clk new_AGEMA_reg_buffer_12450 ( .C (clk), .D (new_AGEMA_signal_25173), .Q (new_AGEMA_signal_25174) ) ;
    buf_clk new_AGEMA_reg_buffer_12453 ( .C (clk), .D (new_AGEMA_signal_25176), .Q (new_AGEMA_signal_25177) ) ;
    buf_clk new_AGEMA_reg_buffer_12456 ( .C (clk), .D (new_AGEMA_signal_25179), .Q (new_AGEMA_signal_25180) ) ;
    buf_clk new_AGEMA_reg_buffer_12459 ( .C (clk), .D (new_AGEMA_signal_25182), .Q (new_AGEMA_signal_25183) ) ;
    buf_clk new_AGEMA_reg_buffer_12462 ( .C (clk), .D (new_AGEMA_signal_25185), .Q (new_AGEMA_signal_25186) ) ;
    buf_clk new_AGEMA_reg_buffer_12465 ( .C (clk), .D (new_AGEMA_signal_25188), .Q (new_AGEMA_signal_25189) ) ;
    buf_clk new_AGEMA_reg_buffer_12468 ( .C (clk), .D (new_AGEMA_signal_25191), .Q (new_AGEMA_signal_25192) ) ;
    buf_clk new_AGEMA_reg_buffer_12471 ( .C (clk), .D (new_AGEMA_signal_25194), .Q (new_AGEMA_signal_25195) ) ;
    buf_clk new_AGEMA_reg_buffer_12474 ( .C (clk), .D (new_AGEMA_signal_25197), .Q (new_AGEMA_signal_25198) ) ;
    buf_clk new_AGEMA_reg_buffer_12477 ( .C (clk), .D (new_AGEMA_signal_25200), .Q (new_AGEMA_signal_25201) ) ;
    buf_clk new_AGEMA_reg_buffer_12480 ( .C (clk), .D (new_AGEMA_signal_25203), .Q (new_AGEMA_signal_25204) ) ;
    buf_clk new_AGEMA_reg_buffer_12483 ( .C (clk), .D (new_AGEMA_signal_25206), .Q (new_AGEMA_signal_25207) ) ;
    buf_clk new_AGEMA_reg_buffer_12486 ( .C (clk), .D (new_AGEMA_signal_25209), .Q (new_AGEMA_signal_25210) ) ;
    buf_clk new_AGEMA_reg_buffer_12489 ( .C (clk), .D (new_AGEMA_signal_25212), .Q (new_AGEMA_signal_25213) ) ;
    buf_clk new_AGEMA_reg_buffer_12492 ( .C (clk), .D (new_AGEMA_signal_25215), .Q (new_AGEMA_signal_25216) ) ;
    buf_clk new_AGEMA_reg_buffer_12495 ( .C (clk), .D (new_AGEMA_signal_25218), .Q (new_AGEMA_signal_25219) ) ;
    buf_clk new_AGEMA_reg_buffer_12498 ( .C (clk), .D (new_AGEMA_signal_25221), .Q (new_AGEMA_signal_25222) ) ;
    buf_clk new_AGEMA_reg_buffer_12501 ( .C (clk), .D (new_AGEMA_signal_25224), .Q (new_AGEMA_signal_25225) ) ;
    buf_clk new_AGEMA_reg_buffer_12504 ( .C (clk), .D (new_AGEMA_signal_25227), .Q (new_AGEMA_signal_25228) ) ;
    buf_clk new_AGEMA_reg_buffer_12507 ( .C (clk), .D (new_AGEMA_signal_25230), .Q (new_AGEMA_signal_25231) ) ;
    buf_clk new_AGEMA_reg_buffer_12510 ( .C (clk), .D (new_AGEMA_signal_25233), .Q (new_AGEMA_signal_25234) ) ;
    buf_clk new_AGEMA_reg_buffer_12513 ( .C (clk), .D (new_AGEMA_signal_25236), .Q (new_AGEMA_signal_25237) ) ;
    buf_clk new_AGEMA_reg_buffer_12516 ( .C (clk), .D (new_AGEMA_signal_25239), .Q (new_AGEMA_signal_25240) ) ;
    buf_clk new_AGEMA_reg_buffer_12519 ( .C (clk), .D (new_AGEMA_signal_25242), .Q (new_AGEMA_signal_25243) ) ;
    buf_clk new_AGEMA_reg_buffer_12522 ( .C (clk), .D (new_AGEMA_signal_25245), .Q (new_AGEMA_signal_25246) ) ;
    buf_clk new_AGEMA_reg_buffer_12525 ( .C (clk), .D (new_AGEMA_signal_25248), .Q (new_AGEMA_signal_25249) ) ;
    buf_clk new_AGEMA_reg_buffer_12528 ( .C (clk), .D (new_AGEMA_signal_25251), .Q (new_AGEMA_signal_25252) ) ;
    buf_clk new_AGEMA_reg_buffer_12531 ( .C (clk), .D (new_AGEMA_signal_25254), .Q (new_AGEMA_signal_25255) ) ;
    buf_clk new_AGEMA_reg_buffer_12534 ( .C (clk), .D (new_AGEMA_signal_25257), .Q (new_AGEMA_signal_25258) ) ;
    buf_clk new_AGEMA_reg_buffer_12537 ( .C (clk), .D (new_AGEMA_signal_25260), .Q (new_AGEMA_signal_25261) ) ;
    buf_clk new_AGEMA_reg_buffer_12540 ( .C (clk), .D (new_AGEMA_signal_25263), .Q (new_AGEMA_signal_25264) ) ;
    buf_clk new_AGEMA_reg_buffer_12543 ( .C (clk), .D (new_AGEMA_signal_25266), .Q (new_AGEMA_signal_25267) ) ;
    buf_clk new_AGEMA_reg_buffer_12546 ( .C (clk), .D (new_AGEMA_signal_25269), .Q (new_AGEMA_signal_25270) ) ;
    buf_clk new_AGEMA_reg_buffer_12549 ( .C (clk), .D (new_AGEMA_signal_25272), .Q (new_AGEMA_signal_25273) ) ;
    buf_clk new_AGEMA_reg_buffer_12552 ( .C (clk), .D (new_AGEMA_signal_25275), .Q (new_AGEMA_signal_25276) ) ;
    buf_clk new_AGEMA_reg_buffer_12555 ( .C (clk), .D (new_AGEMA_signal_25278), .Q (new_AGEMA_signal_25279) ) ;
    buf_clk new_AGEMA_reg_buffer_12558 ( .C (clk), .D (new_AGEMA_signal_25281), .Q (new_AGEMA_signal_25282) ) ;
    buf_clk new_AGEMA_reg_buffer_12561 ( .C (clk), .D (new_AGEMA_signal_25284), .Q (new_AGEMA_signal_25285) ) ;
    buf_clk new_AGEMA_reg_buffer_12564 ( .C (clk), .D (new_AGEMA_signal_25287), .Q (new_AGEMA_signal_25288) ) ;
    buf_clk new_AGEMA_reg_buffer_12567 ( .C (clk), .D (new_AGEMA_signal_25290), .Q (new_AGEMA_signal_25291) ) ;
    buf_clk new_AGEMA_reg_buffer_12570 ( .C (clk), .D (new_AGEMA_signal_25293), .Q (new_AGEMA_signal_25294) ) ;
    buf_clk new_AGEMA_reg_buffer_12573 ( .C (clk), .D (new_AGEMA_signal_25296), .Q (new_AGEMA_signal_25297) ) ;
    buf_clk new_AGEMA_reg_buffer_12576 ( .C (clk), .D (new_AGEMA_signal_25299), .Q (new_AGEMA_signal_25300) ) ;
    buf_clk new_AGEMA_reg_buffer_12579 ( .C (clk), .D (new_AGEMA_signal_25302), .Q (new_AGEMA_signal_25303) ) ;
    buf_clk new_AGEMA_reg_buffer_12582 ( .C (clk), .D (new_AGEMA_signal_25305), .Q (new_AGEMA_signal_25306) ) ;
    buf_clk new_AGEMA_reg_buffer_12585 ( .C (clk), .D (new_AGEMA_signal_25308), .Q (new_AGEMA_signal_25309) ) ;
    buf_clk new_AGEMA_reg_buffer_12588 ( .C (clk), .D (new_AGEMA_signal_25311), .Q (new_AGEMA_signal_25312) ) ;
    buf_clk new_AGEMA_reg_buffer_12591 ( .C (clk), .D (new_AGEMA_signal_25314), .Q (new_AGEMA_signal_25315) ) ;
    buf_clk new_AGEMA_reg_buffer_12594 ( .C (clk), .D (new_AGEMA_signal_25317), .Q (new_AGEMA_signal_25318) ) ;
    buf_clk new_AGEMA_reg_buffer_12597 ( .C (clk), .D (new_AGEMA_signal_25320), .Q (new_AGEMA_signal_25321) ) ;
    buf_clk new_AGEMA_reg_buffer_12600 ( .C (clk), .D (new_AGEMA_signal_25323), .Q (new_AGEMA_signal_25324) ) ;
    buf_clk new_AGEMA_reg_buffer_12603 ( .C (clk), .D (new_AGEMA_signal_25326), .Q (new_AGEMA_signal_25327) ) ;
    buf_clk new_AGEMA_reg_buffer_12606 ( .C (clk), .D (new_AGEMA_signal_25329), .Q (new_AGEMA_signal_25330) ) ;
    buf_clk new_AGEMA_reg_buffer_12609 ( .C (clk), .D (new_AGEMA_signal_25332), .Q (new_AGEMA_signal_25333) ) ;
    buf_clk new_AGEMA_reg_buffer_12612 ( .C (clk), .D (new_AGEMA_signal_25335), .Q (new_AGEMA_signal_25336) ) ;
    buf_clk new_AGEMA_reg_buffer_12615 ( .C (clk), .D (new_AGEMA_signal_25338), .Q (new_AGEMA_signal_25339) ) ;
    buf_clk new_AGEMA_reg_buffer_12618 ( .C (clk), .D (new_AGEMA_signal_25341), .Q (new_AGEMA_signal_25342) ) ;
    buf_clk new_AGEMA_reg_buffer_12621 ( .C (clk), .D (new_AGEMA_signal_25344), .Q (new_AGEMA_signal_25345) ) ;
    buf_clk new_AGEMA_reg_buffer_12624 ( .C (clk), .D (new_AGEMA_signal_25347), .Q (new_AGEMA_signal_25348) ) ;
    buf_clk new_AGEMA_reg_buffer_12627 ( .C (clk), .D (new_AGEMA_signal_25350), .Q (new_AGEMA_signal_25351) ) ;
    buf_clk new_AGEMA_reg_buffer_12630 ( .C (clk), .D (new_AGEMA_signal_25353), .Q (new_AGEMA_signal_25354) ) ;
    buf_clk new_AGEMA_reg_buffer_12633 ( .C (clk), .D (new_AGEMA_signal_25356), .Q (new_AGEMA_signal_25357) ) ;
    buf_clk new_AGEMA_reg_buffer_12636 ( .C (clk), .D (new_AGEMA_signal_25359), .Q (new_AGEMA_signal_25360) ) ;
    buf_clk new_AGEMA_reg_buffer_12639 ( .C (clk), .D (new_AGEMA_signal_25362), .Q (new_AGEMA_signal_25363) ) ;
    buf_clk new_AGEMA_reg_buffer_12642 ( .C (clk), .D (new_AGEMA_signal_25365), .Q (new_AGEMA_signal_25366) ) ;
    buf_clk new_AGEMA_reg_buffer_12645 ( .C (clk), .D (new_AGEMA_signal_25368), .Q (new_AGEMA_signal_25369) ) ;
    buf_clk new_AGEMA_reg_buffer_12648 ( .C (clk), .D (new_AGEMA_signal_25371), .Q (new_AGEMA_signal_25372) ) ;
    buf_clk new_AGEMA_reg_buffer_12651 ( .C (clk), .D (new_AGEMA_signal_25374), .Q (new_AGEMA_signal_25375) ) ;
    buf_clk new_AGEMA_reg_buffer_12654 ( .C (clk), .D (new_AGEMA_signal_25377), .Q (new_AGEMA_signal_25378) ) ;
    buf_clk new_AGEMA_reg_buffer_12657 ( .C (clk), .D (new_AGEMA_signal_25380), .Q (new_AGEMA_signal_25381) ) ;
    buf_clk new_AGEMA_reg_buffer_12660 ( .C (clk), .D (new_AGEMA_signal_25383), .Q (new_AGEMA_signal_25384) ) ;
    buf_clk new_AGEMA_reg_buffer_12663 ( .C (clk), .D (new_AGEMA_signal_25386), .Q (new_AGEMA_signal_25387) ) ;
    buf_clk new_AGEMA_reg_buffer_12666 ( .C (clk), .D (new_AGEMA_signal_25389), .Q (new_AGEMA_signal_25390) ) ;
    buf_clk new_AGEMA_reg_buffer_12669 ( .C (clk), .D (new_AGEMA_signal_25392), .Q (new_AGEMA_signal_25393) ) ;
    buf_clk new_AGEMA_reg_buffer_12672 ( .C (clk), .D (new_AGEMA_signal_25395), .Q (new_AGEMA_signal_25396) ) ;
    buf_clk new_AGEMA_reg_buffer_12675 ( .C (clk), .D (new_AGEMA_signal_25398), .Q (new_AGEMA_signal_25399) ) ;
    buf_clk new_AGEMA_reg_buffer_12678 ( .C (clk), .D (new_AGEMA_signal_25401), .Q (new_AGEMA_signal_25402) ) ;
    buf_clk new_AGEMA_reg_buffer_12681 ( .C (clk), .D (new_AGEMA_signal_25404), .Q (new_AGEMA_signal_25405) ) ;
    buf_clk new_AGEMA_reg_buffer_12684 ( .C (clk), .D (new_AGEMA_signal_25407), .Q (new_AGEMA_signal_25408) ) ;
    buf_clk new_AGEMA_reg_buffer_12687 ( .C (clk), .D (new_AGEMA_signal_25410), .Q (new_AGEMA_signal_25411) ) ;
    buf_clk new_AGEMA_reg_buffer_12690 ( .C (clk), .D (new_AGEMA_signal_25413), .Q (new_AGEMA_signal_25414) ) ;
    buf_clk new_AGEMA_reg_buffer_12693 ( .C (clk), .D (new_AGEMA_signal_25416), .Q (new_AGEMA_signal_25417) ) ;
    buf_clk new_AGEMA_reg_buffer_12696 ( .C (clk), .D (new_AGEMA_signal_25419), .Q (new_AGEMA_signal_25420) ) ;
    buf_clk new_AGEMA_reg_buffer_12699 ( .C (clk), .D (new_AGEMA_signal_25422), .Q (new_AGEMA_signal_25423) ) ;
    buf_clk new_AGEMA_reg_buffer_12702 ( .C (clk), .D (new_AGEMA_signal_25425), .Q (new_AGEMA_signal_25426) ) ;
    buf_clk new_AGEMA_reg_buffer_12705 ( .C (clk), .D (new_AGEMA_signal_25428), .Q (new_AGEMA_signal_25429) ) ;
    buf_clk new_AGEMA_reg_buffer_12708 ( .C (clk), .D (new_AGEMA_signal_25431), .Q (new_AGEMA_signal_25432) ) ;
    buf_clk new_AGEMA_reg_buffer_12711 ( .C (clk), .D (new_AGEMA_signal_25434), .Q (new_AGEMA_signal_25435) ) ;
    buf_clk new_AGEMA_reg_buffer_12714 ( .C (clk), .D (new_AGEMA_signal_25437), .Q (new_AGEMA_signal_25438) ) ;
    buf_clk new_AGEMA_reg_buffer_12717 ( .C (clk), .D (new_AGEMA_signal_25440), .Q (new_AGEMA_signal_25441) ) ;
    buf_clk new_AGEMA_reg_buffer_12720 ( .C (clk), .D (new_AGEMA_signal_25443), .Q (new_AGEMA_signal_25444) ) ;
    buf_clk new_AGEMA_reg_buffer_12723 ( .C (clk), .D (new_AGEMA_signal_25446), .Q (new_AGEMA_signal_25447) ) ;
    buf_clk new_AGEMA_reg_buffer_12726 ( .C (clk), .D (new_AGEMA_signal_25449), .Q (new_AGEMA_signal_25450) ) ;
    buf_clk new_AGEMA_reg_buffer_12729 ( .C (clk), .D (new_AGEMA_signal_25452), .Q (new_AGEMA_signal_25453) ) ;
    buf_clk new_AGEMA_reg_buffer_12732 ( .C (clk), .D (new_AGEMA_signal_25455), .Q (new_AGEMA_signal_25456) ) ;
    buf_clk new_AGEMA_reg_buffer_12735 ( .C (clk), .D (new_AGEMA_signal_25458), .Q (new_AGEMA_signal_25459) ) ;
    buf_clk new_AGEMA_reg_buffer_12738 ( .C (clk), .D (new_AGEMA_signal_25461), .Q (new_AGEMA_signal_25462) ) ;
    buf_clk new_AGEMA_reg_buffer_12741 ( .C (clk), .D (new_AGEMA_signal_25464), .Q (new_AGEMA_signal_25465) ) ;
    buf_clk new_AGEMA_reg_buffer_12744 ( .C (clk), .D (new_AGEMA_signal_25467), .Q (new_AGEMA_signal_25468) ) ;
    buf_clk new_AGEMA_reg_buffer_12747 ( .C (clk), .D (new_AGEMA_signal_25470), .Q (new_AGEMA_signal_25471) ) ;
    buf_clk new_AGEMA_reg_buffer_12750 ( .C (clk), .D (new_AGEMA_signal_25473), .Q (new_AGEMA_signal_25474) ) ;
    buf_clk new_AGEMA_reg_buffer_12753 ( .C (clk), .D (new_AGEMA_signal_25476), .Q (new_AGEMA_signal_25477) ) ;
    buf_clk new_AGEMA_reg_buffer_12756 ( .C (clk), .D (new_AGEMA_signal_25479), .Q (new_AGEMA_signal_25480) ) ;
    buf_clk new_AGEMA_reg_buffer_12759 ( .C (clk), .D (new_AGEMA_signal_25482), .Q (new_AGEMA_signal_25483) ) ;
    buf_clk new_AGEMA_reg_buffer_12762 ( .C (clk), .D (new_AGEMA_signal_25485), .Q (new_AGEMA_signal_25486) ) ;
    buf_clk new_AGEMA_reg_buffer_12765 ( .C (clk), .D (new_AGEMA_signal_25488), .Q (new_AGEMA_signal_25489) ) ;
    buf_clk new_AGEMA_reg_buffer_12768 ( .C (clk), .D (new_AGEMA_signal_25491), .Q (new_AGEMA_signal_25492) ) ;
    buf_clk new_AGEMA_reg_buffer_12771 ( .C (clk), .D (new_AGEMA_signal_25494), .Q (new_AGEMA_signal_25495) ) ;
    buf_clk new_AGEMA_reg_buffer_12774 ( .C (clk), .D (new_AGEMA_signal_25497), .Q (new_AGEMA_signal_25498) ) ;
    buf_clk new_AGEMA_reg_buffer_12777 ( .C (clk), .D (new_AGEMA_signal_25500), .Q (new_AGEMA_signal_25501) ) ;
    buf_clk new_AGEMA_reg_buffer_12780 ( .C (clk), .D (new_AGEMA_signal_25503), .Q (new_AGEMA_signal_25504) ) ;
    buf_clk new_AGEMA_reg_buffer_12783 ( .C (clk), .D (new_AGEMA_signal_25506), .Q (new_AGEMA_signal_25507) ) ;
    buf_clk new_AGEMA_reg_buffer_12786 ( .C (clk), .D (new_AGEMA_signal_25509), .Q (new_AGEMA_signal_25510) ) ;
    buf_clk new_AGEMA_reg_buffer_12789 ( .C (clk), .D (new_AGEMA_signal_25512), .Q (new_AGEMA_signal_25513) ) ;
    buf_clk new_AGEMA_reg_buffer_12792 ( .C (clk), .D (new_AGEMA_signal_25515), .Q (new_AGEMA_signal_25516) ) ;
    buf_clk new_AGEMA_reg_buffer_12795 ( .C (clk), .D (new_AGEMA_signal_25518), .Q (new_AGEMA_signal_25519) ) ;
    buf_clk new_AGEMA_reg_buffer_12798 ( .C (clk), .D (new_AGEMA_signal_25521), .Q (new_AGEMA_signal_25522) ) ;
    buf_clk new_AGEMA_reg_buffer_12801 ( .C (clk), .D (new_AGEMA_signal_25524), .Q (new_AGEMA_signal_25525) ) ;
    buf_clk new_AGEMA_reg_buffer_12804 ( .C (clk), .D (new_AGEMA_signal_25527), .Q (new_AGEMA_signal_25528) ) ;
    buf_clk new_AGEMA_reg_buffer_12807 ( .C (clk), .D (new_AGEMA_signal_25530), .Q (new_AGEMA_signal_25531) ) ;
    buf_clk new_AGEMA_reg_buffer_12811 ( .C (clk), .D (new_AGEMA_signal_25534), .Q (new_AGEMA_signal_25535) ) ;
    buf_clk new_AGEMA_reg_buffer_12815 ( .C (clk), .D (new_AGEMA_signal_25538), .Q (new_AGEMA_signal_25539) ) ;
    buf_clk new_AGEMA_reg_buffer_12819 ( .C (clk), .D (new_AGEMA_signal_25542), .Q (new_AGEMA_signal_25543) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(2), .pipeline(1)) U858 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .a ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U859 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_12218, new_AGEMA_signal_12217, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U860 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_11834, new_AGEMA_signal_11833, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U861 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_11396, new_AGEMA_signal_11395, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U862 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U863 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_11840, new_AGEMA_signal_11839, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U864 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U865 ( .s (new_AGEMA_signal_17656), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .a ({new_AGEMA_signal_11450, new_AGEMA_signal_11449, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U866 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .a ({new_AGEMA_signal_12014, new_AGEMA_signal_12013, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U867 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_12224, new_AGEMA_signal_12223, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U868 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_11444, new_AGEMA_signal_11443, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U869 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .a ({new_AGEMA_signal_11642, new_AGEMA_signal_11641, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_11846, new_AGEMA_signal_11845, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U870 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U871 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U872 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .a ({new_AGEMA_signal_11438, new_AGEMA_signal_11437, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_11852, new_AGEMA_signal_11851, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U873 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U874 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .a ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U875 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .a ({new_AGEMA_signal_12008, new_AGEMA_signal_12007, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U876 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_12230, new_AGEMA_signal_12229, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U877 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_11426, new_AGEMA_signal_11425, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U878 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_11858, new_AGEMA_signal_11857, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U879 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U880 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .a ({new_AGEMA_signal_12086, new_AGEMA_signal_12085, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U881 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .a ({new_AGEMA_signal_11420, new_AGEMA_signal_11419, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U882 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_12002, new_AGEMA_signal_12001, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U883 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .a ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_11864, new_AGEMA_signal_11863, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U884 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .a ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_12236, new_AGEMA_signal_12235, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U885 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U886 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U887 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U888 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_11870, new_AGEMA_signal_11869, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U889 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U890 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_11636, new_AGEMA_signal_11635, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U891 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U892 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_11876, new_AGEMA_signal_11875, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U893 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .a ({new_AGEMA_signal_11630, new_AGEMA_signal_11629, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U894 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_12242, new_AGEMA_signal_12241, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U895 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .a ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U896 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .a ({new_AGEMA_signal_12080, new_AGEMA_signal_12079, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U897 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U898 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_12248, new_AGEMA_signal_12247, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U899 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_11618, new_AGEMA_signal_11617, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_11882, new_AGEMA_signal_11881, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U900 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U901 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U902 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .a ({new_AGEMA_signal_11612, new_AGEMA_signal_11611, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_11888, new_AGEMA_signal_11887, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U903 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_12074, new_AGEMA_signal_12073, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U904 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .a ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U905 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .a ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U906 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_12254, new_AGEMA_signal_12253, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U907 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U908 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .a ({new_AGEMA_signal_11600, new_AGEMA_signal_11599, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_11894, new_AGEMA_signal_11893, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U909 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U910 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U911 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .a ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_11900, new_AGEMA_signal_11899, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U912 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U913 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .a ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U914 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .a ({new_AGEMA_signal_12044, new_AGEMA_signal_12043, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U915 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_12260, new_AGEMA_signal_12259, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U916 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U917 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_11906, new_AGEMA_signal_11905, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U918 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_11522, new_AGEMA_signal_11521, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U919 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .a ({new_AGEMA_signal_12068, new_AGEMA_signal_12067, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U920 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .a ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U921 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U922 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .a ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_11912, new_AGEMA_signal_11911, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U923 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .a ({new_AGEMA_signal_12062, new_AGEMA_signal_12061, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_12266, new_AGEMA_signal_12265, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U924 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U925 ( .s (new_AGEMA_signal_17680), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U926 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_11570, new_AGEMA_signal_11569, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U927 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_11918, new_AGEMA_signal_11917, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U928 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .a ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U929 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U930 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_12272, new_AGEMA_signal_12271, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U931 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .a ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U932 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .a ({new_AGEMA_signal_12056, new_AGEMA_signal_12055, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U933 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U934 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_11924, new_AGEMA_signal_11923, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U935 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_11552, new_AGEMA_signal_11551, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U936 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U937 ( .s (new_AGEMA_signal_17676), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .a ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_11930, new_AGEMA_signal_11929, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U938 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_12050, new_AGEMA_signal_12049, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_12278, new_AGEMA_signal_12277, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U939 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .a ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U940 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U941 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U942 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U943 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_11936, new_AGEMA_signal_11935, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U944 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_11534, new_AGEMA_signal_11533, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U945 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U946 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .a ({new_AGEMA_signal_11516, new_AGEMA_signal_11515, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_11942, new_AGEMA_signal_11941, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U947 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_12284, new_AGEMA_signal_12283, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U948 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .a ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U949 ( .s (new_AGEMA_signal_17672), .b ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .a ({new_AGEMA_signal_12020, new_AGEMA_signal_12019, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U950 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U951 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_11462, new_AGEMA_signal_11461, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U952 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_11588, new_AGEMA_signal_11587, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_11948, new_AGEMA_signal_11947, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U953 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U954 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U955 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .a ({new_AGEMA_signal_11456, new_AGEMA_signal_11455, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_11954, new_AGEMA_signal_11953, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U956 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_12290, new_AGEMA_signal_12289, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U957 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .a ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U958 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .a ({new_AGEMA_signal_12038, new_AGEMA_signal_12037, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U959 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U960 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U961 ( .s (new_AGEMA_signal_17668), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_11960, new_AGEMA_signal_11959, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U962 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_11504, new_AGEMA_signal_11503, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U963 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U964 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .a ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_11966, new_AGEMA_signal_11965, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U965 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_12296, new_AGEMA_signal_12295, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U966 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .a ({new_AGEMA_signal_11498, new_AGEMA_signal_11497, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U967 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .a ({new_AGEMA_signal_12032, new_AGEMA_signal_12031, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U968 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U969 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U970 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_11972, new_AGEMA_signal_11971, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U971 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_11486, new_AGEMA_signal_11485, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U972 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .a ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U973 ( .s (new_AGEMA_signal_17664), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_12026, new_AGEMA_signal_12025, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_12302, new_AGEMA_signal_12301, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U974 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .a ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_11978, new_AGEMA_signal_11977, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U975 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .a ({new_AGEMA_signal_11480, new_AGEMA_signal_11479, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U976 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .a ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U977 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U978 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_11474, new_AGEMA_signal_11473, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U979 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_11984, new_AGEMA_signal_11983, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U980 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_11468, new_AGEMA_signal_11467, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U981 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .a ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U982 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_12308, new_AGEMA_signal_12307, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U983 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .a ({new_AGEMA_signal_11408, new_AGEMA_signal_11407, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_11990, new_AGEMA_signal_11989, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U984 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .a ({new_AGEMA_signal_11996, new_AGEMA_signal_11995, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) U985 ( .s (new_AGEMA_signal_17660), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, RoundOutput[0]}), .a ({new_AGEMA_signal_17696, new_AGEMA_signal_17692, new_AGEMA_signal_17688}), .c ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, RoundOutput[1]}), .a ({new_AGEMA_signal_17708, new_AGEMA_signal_17704, new_AGEMA_signal_17700}), .c ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11894, new_AGEMA_signal_11893, RoundOutput[2]}), .a ({new_AGEMA_signal_17720, new_AGEMA_signal_17716, new_AGEMA_signal_17712}), .c ({new_AGEMA_signal_12320, new_AGEMA_signal_12319, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, RoundOutput[3]}), .a ({new_AGEMA_signal_17732, new_AGEMA_signal_17728, new_AGEMA_signal_17724}), .c ({new_AGEMA_signal_12668, new_AGEMA_signal_12667, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12272, new_AGEMA_signal_12271, RoundOutput[4]}), .a ({new_AGEMA_signal_17744, new_AGEMA_signal_17740, new_AGEMA_signal_17736}), .c ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, RoundOutput[5]}), .a ({new_AGEMA_signal_17756, new_AGEMA_signal_17752, new_AGEMA_signal_17748}), .c ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11948, new_AGEMA_signal_11947, RoundOutput[6]}), .a ({new_AGEMA_signal_17768, new_AGEMA_signal_17764, new_AGEMA_signal_17760}), .c ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, RoundOutput[7]}), .a ({new_AGEMA_signal_17780, new_AGEMA_signal_17776, new_AGEMA_signal_17772}), .c ({new_AGEMA_signal_12332, new_AGEMA_signal_12331, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11978, new_AGEMA_signal_11977, RoundOutput[8]}), .a ({new_AGEMA_signal_17792, new_AGEMA_signal_17788, new_AGEMA_signal_17784}), .c ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, RoundOutput[9]}), .a ({new_AGEMA_signal_17804, new_AGEMA_signal_17800, new_AGEMA_signal_17796}), .c ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11846, new_AGEMA_signal_11845, RoundOutput[10]}), .a ({new_AGEMA_signal_17816, new_AGEMA_signal_17812, new_AGEMA_signal_17808}), .c ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, RoundOutput[11]}), .a ({new_AGEMA_signal_17828, new_AGEMA_signal_17824, new_AGEMA_signal_17820}), .c ({new_AGEMA_signal_12680, new_AGEMA_signal_12679, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, RoundOutput[12]}), .a ({new_AGEMA_signal_17840, new_AGEMA_signal_17836, new_AGEMA_signal_17832}), .c ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, RoundOutput[13]}), .a ({new_AGEMA_signal_17852, new_AGEMA_signal_17848, new_AGEMA_signal_17844}), .c ({new_AGEMA_signal_12344, new_AGEMA_signal_12343, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, RoundOutput[14]}), .a ({new_AGEMA_signal_17864, new_AGEMA_signal_17860, new_AGEMA_signal_17856}), .c ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11876, new_AGEMA_signal_11875, RoundOutput[15]}), .a ({new_AGEMA_signal_17876, new_AGEMA_signal_17872, new_AGEMA_signal_17868}), .c ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, RoundOutput[16]}), .a ({new_AGEMA_signal_17888, new_AGEMA_signal_17884, new_AGEMA_signal_17880}), .c ({new_AGEMA_signal_12356, new_AGEMA_signal_12355, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12242, new_AGEMA_signal_12241, RoundOutput[17]}), .a ({new_AGEMA_signal_17900, new_AGEMA_signal_17896, new_AGEMA_signal_17892}), .c ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, RoundOutput[18]}), .a ({new_AGEMA_signal_17912, new_AGEMA_signal_17908, new_AGEMA_signal_17904}), .c ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, RoundOutput[19]}), .a ({new_AGEMA_signal_17924, new_AGEMA_signal_17920, new_AGEMA_signal_17916}), .c ({new_AGEMA_signal_12692, new_AGEMA_signal_12691, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12248, new_AGEMA_signal_12247, RoundOutput[20]}), .a ({new_AGEMA_signal_17936, new_AGEMA_signal_17932, new_AGEMA_signal_17928}), .c ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11882, new_AGEMA_signal_11881, RoundOutput[21]}), .a ({new_AGEMA_signal_17948, new_AGEMA_signal_17944, new_AGEMA_signal_17940}), .c ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, RoundOutput[22]}), .a ({new_AGEMA_signal_17960, new_AGEMA_signal_17956, new_AGEMA_signal_17952}), .c ({new_AGEMA_signal_12368, new_AGEMA_signal_12367, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, RoundOutput[23]}), .a ({new_AGEMA_signal_17972, new_AGEMA_signal_17968, new_AGEMA_signal_17964}), .c ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11888, new_AGEMA_signal_11887, RoundOutput[24]}), .a ({new_AGEMA_signal_17984, new_AGEMA_signal_17980, new_AGEMA_signal_17976}), .c ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, RoundOutput[25]}), .a ({new_AGEMA_signal_17996, new_AGEMA_signal_17992, new_AGEMA_signal_17988}), .c ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, RoundOutput[26]}), .a ({new_AGEMA_signal_18008, new_AGEMA_signal_18004, new_AGEMA_signal_18000}), .c ({new_AGEMA_signal_12380, new_AGEMA_signal_12379, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, RoundOutput[27]}), .a ({new_AGEMA_signal_18020, new_AGEMA_signal_18016, new_AGEMA_signal_18012}), .c ({new_AGEMA_signal_12704, new_AGEMA_signal_12703, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12254, new_AGEMA_signal_12253, RoundOutput[28]}), .a ({new_AGEMA_signal_18032, new_AGEMA_signal_18028, new_AGEMA_signal_18024}), .c ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, RoundOutput[29]}), .a ({new_AGEMA_signal_18044, new_AGEMA_signal_18040, new_AGEMA_signal_18036}), .c ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, RoundOutput[30]}), .a ({new_AGEMA_signal_18056, new_AGEMA_signal_18052, new_AGEMA_signal_18048}), .c ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, RoundOutput[31]}), .a ({new_AGEMA_signal_18068, new_AGEMA_signal_18064, new_AGEMA_signal_18060}), .c ({new_AGEMA_signal_12392, new_AGEMA_signal_12391, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11900, new_AGEMA_signal_11899, RoundOutput[32]}), .a ({new_AGEMA_signal_18080, new_AGEMA_signal_18076, new_AGEMA_signal_18072}), .c ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, RoundOutput[33]}), .a ({new_AGEMA_signal_18092, new_AGEMA_signal_18088, new_AGEMA_signal_18084}), .c ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, RoundOutput[34]}), .a ({new_AGEMA_signal_18104, new_AGEMA_signal_18100, new_AGEMA_signal_18096}), .c ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, RoundOutput[35]}), .a ({new_AGEMA_signal_18116, new_AGEMA_signal_18112, new_AGEMA_signal_18108}), .c ({new_AGEMA_signal_12716, new_AGEMA_signal_12715, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12260, new_AGEMA_signal_12259, RoundOutput[36]}), .a ({new_AGEMA_signal_18128, new_AGEMA_signal_18124, new_AGEMA_signal_18120}), .c ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, RoundOutput[37]}), .a ({new_AGEMA_signal_18140, new_AGEMA_signal_18136, new_AGEMA_signal_18132}), .c ({new_AGEMA_signal_12404, new_AGEMA_signal_12403, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11906, new_AGEMA_signal_11905, RoundOutput[38]}), .a ({new_AGEMA_signal_18152, new_AGEMA_signal_18148, new_AGEMA_signal_18144}), .c ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, RoundOutput[39]}), .a ({new_AGEMA_signal_18164, new_AGEMA_signal_18160, new_AGEMA_signal_18156}), .c ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, RoundOutput[40]}), .a ({new_AGEMA_signal_18176, new_AGEMA_signal_18172, new_AGEMA_signal_18168}), .c ({new_AGEMA_signal_12416, new_AGEMA_signal_12415, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, RoundOutput[41]}), .a ({new_AGEMA_signal_18188, new_AGEMA_signal_18184, new_AGEMA_signal_18180}), .c ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11912, new_AGEMA_signal_11911, RoundOutput[42]}), .a ({new_AGEMA_signal_18200, new_AGEMA_signal_18196, new_AGEMA_signal_18192}), .c ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12266, new_AGEMA_signal_12265, RoundOutput[43]}), .a ({new_AGEMA_signal_18212, new_AGEMA_signal_18208, new_AGEMA_signal_18204}), .c ({new_AGEMA_signal_12728, new_AGEMA_signal_12727, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, RoundOutput[44]}), .a ({new_AGEMA_signal_18224, new_AGEMA_signal_18220, new_AGEMA_signal_18216}), .c ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, RoundOutput[45]}), .a ({new_AGEMA_signal_18236, new_AGEMA_signal_18232, new_AGEMA_signal_18228}), .c ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, RoundOutput[46]}), .a ({new_AGEMA_signal_18248, new_AGEMA_signal_18244, new_AGEMA_signal_18240}), .c ({new_AGEMA_signal_12428, new_AGEMA_signal_12427, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11918, new_AGEMA_signal_11917, RoundOutput[47]}), .a ({new_AGEMA_signal_18260, new_AGEMA_signal_18256, new_AGEMA_signal_18252}), .c ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, RoundOutput[48]}), .a ({new_AGEMA_signal_18272, new_AGEMA_signal_18268, new_AGEMA_signal_18264}), .c ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, RoundOutput[49]}), .a ({new_AGEMA_signal_18284, new_AGEMA_signal_18280, new_AGEMA_signal_18276}), .c ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, RoundOutput[50]}), .a ({new_AGEMA_signal_18296, new_AGEMA_signal_18292, new_AGEMA_signal_18288}), .c ({new_AGEMA_signal_12440, new_AGEMA_signal_12439, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, RoundOutput[51]}), .a ({new_AGEMA_signal_18308, new_AGEMA_signal_18304, new_AGEMA_signal_18300}), .c ({new_AGEMA_signal_12740, new_AGEMA_signal_12739, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, RoundOutput[52]}), .a ({new_AGEMA_signal_18320, new_AGEMA_signal_18316, new_AGEMA_signal_18312}), .c ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11924, new_AGEMA_signal_11923, RoundOutput[53]}), .a ({new_AGEMA_signal_18332, new_AGEMA_signal_18328, new_AGEMA_signal_18324}), .c ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, RoundOutput[54]}), .a ({new_AGEMA_signal_18344, new_AGEMA_signal_18340, new_AGEMA_signal_18336}), .c ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, RoundOutput[55]}), .a ({new_AGEMA_signal_18356, new_AGEMA_signal_18352, new_AGEMA_signal_18348}), .c ({new_AGEMA_signal_12452, new_AGEMA_signal_12451, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11930, new_AGEMA_signal_11929, RoundOutput[56]}), .a ({new_AGEMA_signal_18368, new_AGEMA_signal_18364, new_AGEMA_signal_18360}), .c ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12278, new_AGEMA_signal_12277, RoundOutput[57]}), .a ({new_AGEMA_signal_18380, new_AGEMA_signal_18376, new_AGEMA_signal_18372}), .c ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, RoundOutput[58]}), .a ({new_AGEMA_signal_18392, new_AGEMA_signal_18388, new_AGEMA_signal_18384}), .c ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, RoundOutput[59]}), .a ({new_AGEMA_signal_18404, new_AGEMA_signal_18400, new_AGEMA_signal_18396}), .c ({new_AGEMA_signal_12752, new_AGEMA_signal_12751, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, RoundOutput[60]}), .a ({new_AGEMA_signal_18416, new_AGEMA_signal_18412, new_AGEMA_signal_18408}), .c ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11936, new_AGEMA_signal_11935, RoundOutput[61]}), .a ({new_AGEMA_signal_18428, new_AGEMA_signal_18424, new_AGEMA_signal_18420}), .c ({new_AGEMA_signal_12464, new_AGEMA_signal_12463, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, RoundOutput[62]}), .a ({new_AGEMA_signal_18440, new_AGEMA_signal_18436, new_AGEMA_signal_18432}), .c ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, RoundOutput[63]}), .a ({new_AGEMA_signal_18452, new_AGEMA_signal_18448, new_AGEMA_signal_18444}), .c ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11942, new_AGEMA_signal_11941, RoundOutput[64]}), .a ({new_AGEMA_signal_18464, new_AGEMA_signal_18460, new_AGEMA_signal_18456}), .c ({new_AGEMA_signal_12476, new_AGEMA_signal_12475, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12284, new_AGEMA_signal_12283, RoundOutput[65]}), .a ({new_AGEMA_signal_18476, new_AGEMA_signal_18472, new_AGEMA_signal_18468}), .c ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, RoundOutput[66]}), .a ({new_AGEMA_signal_18488, new_AGEMA_signal_18484, new_AGEMA_signal_18480}), .c ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, RoundOutput[67]}), .a ({new_AGEMA_signal_18500, new_AGEMA_signal_18496, new_AGEMA_signal_18492}), .c ({new_AGEMA_signal_12764, new_AGEMA_signal_12763, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, RoundOutput[68]}), .a ({new_AGEMA_signal_18512, new_AGEMA_signal_18508, new_AGEMA_signal_18504}), .c ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, RoundOutput[69]}), .a ({new_AGEMA_signal_18524, new_AGEMA_signal_18520, new_AGEMA_signal_18516}), .c ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, RoundOutput[70]}), .a ({new_AGEMA_signal_18536, new_AGEMA_signal_18532, new_AGEMA_signal_18528}), .c ({new_AGEMA_signal_12488, new_AGEMA_signal_12487, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, RoundOutput[71]}), .a ({new_AGEMA_signal_18548, new_AGEMA_signal_18544, new_AGEMA_signal_18540}), .c ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11954, new_AGEMA_signal_11953, RoundOutput[72]}), .a ({new_AGEMA_signal_18560, new_AGEMA_signal_18556, new_AGEMA_signal_18552}), .c ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12290, new_AGEMA_signal_12289, RoundOutput[73]}), .a ({new_AGEMA_signal_18572, new_AGEMA_signal_18568, new_AGEMA_signal_18564}), .c ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, RoundOutput[74]}), .a ({new_AGEMA_signal_18584, new_AGEMA_signal_18580, new_AGEMA_signal_18576}), .c ({new_AGEMA_signal_12500, new_AGEMA_signal_12499, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, RoundOutput[75]}), .a ({new_AGEMA_signal_18596, new_AGEMA_signal_18592, new_AGEMA_signal_18588}), .c ({new_AGEMA_signal_12776, new_AGEMA_signal_12775, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, RoundOutput[76]}), .a ({new_AGEMA_signal_18608, new_AGEMA_signal_18604, new_AGEMA_signal_18600}), .c ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, RoundOutput[77]}), .a ({new_AGEMA_signal_18620, new_AGEMA_signal_18616, new_AGEMA_signal_18612}), .c ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11960, new_AGEMA_signal_11959, RoundOutput[78]}), .a ({new_AGEMA_signal_18632, new_AGEMA_signal_18628, new_AGEMA_signal_18624}), .c ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, RoundOutput[79]}), .a ({new_AGEMA_signal_18644, new_AGEMA_signal_18640, new_AGEMA_signal_18636}), .c ({new_AGEMA_signal_12512, new_AGEMA_signal_12511, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11966, new_AGEMA_signal_11965, RoundOutput[80]}), .a ({new_AGEMA_signal_18656, new_AGEMA_signal_18652, new_AGEMA_signal_18648}), .c ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12296, new_AGEMA_signal_12295, RoundOutput[81]}), .a ({new_AGEMA_signal_18668, new_AGEMA_signal_18664, new_AGEMA_signal_18660}), .c ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, RoundOutput[82]}), .a ({new_AGEMA_signal_18680, new_AGEMA_signal_18676, new_AGEMA_signal_18672}), .c ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, RoundOutput[83]}), .a ({new_AGEMA_signal_18692, new_AGEMA_signal_18688, new_AGEMA_signal_18684}), .c ({new_AGEMA_signal_12788, new_AGEMA_signal_12787, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, RoundOutput[84]}), .a ({new_AGEMA_signal_18704, new_AGEMA_signal_18700, new_AGEMA_signal_18696}), .c ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, RoundOutput[85]}), .a ({new_AGEMA_signal_18716, new_AGEMA_signal_18712, new_AGEMA_signal_18708}), .c ({new_AGEMA_signal_12524, new_AGEMA_signal_12523, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11972, new_AGEMA_signal_11971, RoundOutput[86]}), .a ({new_AGEMA_signal_18728, new_AGEMA_signal_18724, new_AGEMA_signal_18720}), .c ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, RoundOutput[87]}), .a ({new_AGEMA_signal_18740, new_AGEMA_signal_18736, new_AGEMA_signal_18732}), .c ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, RoundOutput[88]}), .a ({new_AGEMA_signal_18752, new_AGEMA_signal_18748, new_AGEMA_signal_18744}), .c ({new_AGEMA_signal_12536, new_AGEMA_signal_12535, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12302, new_AGEMA_signal_12301, RoundOutput[89]}), .a ({new_AGEMA_signal_18764, new_AGEMA_signal_18760, new_AGEMA_signal_18756}), .c ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, RoundOutput[90]}), .a ({new_AGEMA_signal_18776, new_AGEMA_signal_18772, new_AGEMA_signal_18768}), .c ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, RoundOutput[91]}), .a ({new_AGEMA_signal_18788, new_AGEMA_signal_18784, new_AGEMA_signal_18780}), .c ({new_AGEMA_signal_12800, new_AGEMA_signal_12799, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, RoundOutput[92]}), .a ({new_AGEMA_signal_18800, new_AGEMA_signal_18796, new_AGEMA_signal_18792}), .c ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, RoundOutput[93]}), .a ({new_AGEMA_signal_18812, new_AGEMA_signal_18808, new_AGEMA_signal_18804}), .c ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11984, new_AGEMA_signal_11983, RoundOutput[94]}), .a ({new_AGEMA_signal_18824, new_AGEMA_signal_18820, new_AGEMA_signal_18816}), .c ({new_AGEMA_signal_12548, new_AGEMA_signal_12547, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, RoundOutput[95]}), .a ({new_AGEMA_signal_18836, new_AGEMA_signal_18832, new_AGEMA_signal_18828}), .c ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, RoundOutput[96]}), .a ({new_AGEMA_signal_18848, new_AGEMA_signal_18844, new_AGEMA_signal_18840}), .c ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12308, new_AGEMA_signal_12307, RoundOutput[97]}), .a ({new_AGEMA_signal_18860, new_AGEMA_signal_18856, new_AGEMA_signal_18852}), .c ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11990, new_AGEMA_signal_11989, RoundOutput[98]}), .a ({new_AGEMA_signal_18872, new_AGEMA_signal_18868, new_AGEMA_signal_18864}), .c ({new_AGEMA_signal_12560, new_AGEMA_signal_12559, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, RoundOutput[99]}), .a ({new_AGEMA_signal_18884, new_AGEMA_signal_18880, new_AGEMA_signal_18876}), .c ({new_AGEMA_signal_12812, new_AGEMA_signal_12811, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12218, new_AGEMA_signal_12217, RoundOutput[100]}), .a ({new_AGEMA_signal_18896, new_AGEMA_signal_18892, new_AGEMA_signal_18888}), .c ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11834, new_AGEMA_signal_11833, RoundOutput[101]}), .a ({new_AGEMA_signal_18908, new_AGEMA_signal_18904, new_AGEMA_signal_18900}), .c ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, RoundOutput[102]}), .a ({new_AGEMA_signal_18920, new_AGEMA_signal_18916, new_AGEMA_signal_18912}), .c ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, RoundOutput[103]}), .a ({new_AGEMA_signal_18932, new_AGEMA_signal_18928, new_AGEMA_signal_18924}), .c ({new_AGEMA_signal_12572, new_AGEMA_signal_12571, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11840, new_AGEMA_signal_11839, RoundOutput[104]}), .a ({new_AGEMA_signal_18944, new_AGEMA_signal_18940, new_AGEMA_signal_18936}), .c ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, RoundOutput[105]}), .a ({new_AGEMA_signal_18956, new_AGEMA_signal_18952, new_AGEMA_signal_18948}), .c ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, RoundOutput[106]}), .a ({new_AGEMA_signal_18968, new_AGEMA_signal_18964, new_AGEMA_signal_18960}), .c ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, RoundOutput[107]}), .a ({new_AGEMA_signal_18980, new_AGEMA_signal_18976, new_AGEMA_signal_18972}), .c ({new_AGEMA_signal_12824, new_AGEMA_signal_12823, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12224, new_AGEMA_signal_12223, RoundOutput[108]}), .a ({new_AGEMA_signal_18992, new_AGEMA_signal_18988, new_AGEMA_signal_18984}), .c ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, RoundOutput[109]}), .a ({new_AGEMA_signal_19004, new_AGEMA_signal_19000, new_AGEMA_signal_18996}), .c ({new_AGEMA_signal_12584, new_AGEMA_signal_12583, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, RoundOutput[110]}), .a ({new_AGEMA_signal_19016, new_AGEMA_signal_19012, new_AGEMA_signal_19008}), .c ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, RoundOutput[111]}), .a ({new_AGEMA_signal_19028, new_AGEMA_signal_19024, new_AGEMA_signal_19020}), .c ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11852, new_AGEMA_signal_11851, RoundOutput[112]}), .a ({new_AGEMA_signal_19040, new_AGEMA_signal_19036, new_AGEMA_signal_19032}), .c ({new_AGEMA_signal_12596, new_AGEMA_signal_12595, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, RoundOutput[113]}), .a ({new_AGEMA_signal_19052, new_AGEMA_signal_19048, new_AGEMA_signal_19044}), .c ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, RoundOutput[114]}), .a ({new_AGEMA_signal_19064, new_AGEMA_signal_19060, new_AGEMA_signal_19056}), .c ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, RoundOutput[115]}), .a ({new_AGEMA_signal_19076, new_AGEMA_signal_19072, new_AGEMA_signal_19068}), .c ({new_AGEMA_signal_12836, new_AGEMA_signal_12835, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12230, new_AGEMA_signal_12229, RoundOutput[116]}), .a ({new_AGEMA_signal_19088, new_AGEMA_signal_19084, new_AGEMA_signal_19080}), .c ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, RoundOutput[117]}), .a ({new_AGEMA_signal_19100, new_AGEMA_signal_19096, new_AGEMA_signal_19092}), .c ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11858, new_AGEMA_signal_11857, RoundOutput[118]}), .a ({new_AGEMA_signal_19112, new_AGEMA_signal_19108, new_AGEMA_signal_19104}), .c ({new_AGEMA_signal_12608, new_AGEMA_signal_12607, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, RoundOutput[119]}), .a ({new_AGEMA_signal_19124, new_AGEMA_signal_19120, new_AGEMA_signal_19116}), .c ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, RoundOutput[120]}), .a ({new_AGEMA_signal_19136, new_AGEMA_signal_19132, new_AGEMA_signal_19128}), .c ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, RoundOutput[121]}), .a ({new_AGEMA_signal_19148, new_AGEMA_signal_19144, new_AGEMA_signal_19140}), .c ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11864, new_AGEMA_signal_11863, RoundOutput[122]}), .a ({new_AGEMA_signal_19160, new_AGEMA_signal_19156, new_AGEMA_signal_19152}), .c ({new_AGEMA_signal_12620, new_AGEMA_signal_12619, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12236, new_AGEMA_signal_12235, RoundOutput[123]}), .a ({new_AGEMA_signal_19172, new_AGEMA_signal_19168, new_AGEMA_signal_19164}), .c ({new_AGEMA_signal_12848, new_AGEMA_signal_12847, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, RoundOutput[124]}), .a ({new_AGEMA_signal_19184, new_AGEMA_signal_19180, new_AGEMA_signal_19176}), .c ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, RoundOutput[125]}), .a ({new_AGEMA_signal_19196, new_AGEMA_signal_19192, new_AGEMA_signal_19188}), .c ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, RoundOutput[126]}), .a ({new_AGEMA_signal_19208, new_AGEMA_signal_19204, new_AGEMA_signal_19200}), .c ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11870, new_AGEMA_signal_11869, RoundOutput[127]}), .a ({new_AGEMA_signal_19220, new_AGEMA_signal_19216, new_AGEMA_signal_19212}), .c ({new_AGEMA_signal_12632, new_AGEMA_signal_12631, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_19229, new_AGEMA_signal_19226, new_AGEMA_signal_19223}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_19238, new_AGEMA_signal_19235, new_AGEMA_signal_19232}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_8102, new_AGEMA_signal_8101, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_19247, new_AGEMA_signal_19244, new_AGEMA_signal_19241}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_19256, new_AGEMA_signal_19253, new_AGEMA_signal_19250}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_19265, new_AGEMA_signal_19262, new_AGEMA_signal_19259}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_19274, new_AGEMA_signal_19271, new_AGEMA_signal_19268}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_19283, new_AGEMA_signal_19280, new_AGEMA_signal_19277}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_19292, new_AGEMA_signal_19289, new_AGEMA_signal_19286}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_19301, new_AGEMA_signal_19298, new_AGEMA_signal_19295}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_19310, new_AGEMA_signal_19307, new_AGEMA_signal_19304}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_19319, new_AGEMA_signal_19316, new_AGEMA_signal_19313}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_19328, new_AGEMA_signal_19325, new_AGEMA_signal_19322}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_19337, new_AGEMA_signal_19334, new_AGEMA_signal_19331}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_19346, new_AGEMA_signal_19343, new_AGEMA_signal_19340}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_8114, new_AGEMA_signal_8113, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_19355, new_AGEMA_signal_19352, new_AGEMA_signal_19349}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_19364, new_AGEMA_signal_19361, new_AGEMA_signal_19358}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_19373, new_AGEMA_signal_19370, new_AGEMA_signal_19367}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_19382, new_AGEMA_signal_19379, new_AGEMA_signal_19376}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_8102, new_AGEMA_signal_8101, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_8114, new_AGEMA_signal_8113, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_8108, new_AGEMA_signal_8107, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9806, new_AGEMA_signal_9805, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_9812, new_AGEMA_signal_9811, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9818, new_AGEMA_signal_9817, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_9824, new_AGEMA_signal_9823, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_9818, new_AGEMA_signal_9817, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9812, new_AGEMA_signal_9811, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_9824, new_AGEMA_signal_9823, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_9806, new_AGEMA_signal_9805, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_19391, new_AGEMA_signal_19388, new_AGEMA_signal_19385}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_19400, new_AGEMA_signal_19397, new_AGEMA_signal_19394}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_8126, new_AGEMA_signal_8125, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_19409, new_AGEMA_signal_19406, new_AGEMA_signal_19403}), .clk (clk), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_19418, new_AGEMA_signal_19415, new_AGEMA_signal_19412}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_19427, new_AGEMA_signal_19424, new_AGEMA_signal_19421}), .clk (clk), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_19436, new_AGEMA_signal_19433, new_AGEMA_signal_19430}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_19445, new_AGEMA_signal_19442, new_AGEMA_signal_19439}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_19454, new_AGEMA_signal_19451, new_AGEMA_signal_19448}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_19463, new_AGEMA_signal_19460, new_AGEMA_signal_19457}), .clk (clk), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_19472, new_AGEMA_signal_19469, new_AGEMA_signal_19466}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_19481, new_AGEMA_signal_19478, new_AGEMA_signal_19475}), .clk (clk), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_19490, new_AGEMA_signal_19487, new_AGEMA_signal_19484}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_19499, new_AGEMA_signal_19496, new_AGEMA_signal_19493}), .clk (clk), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_19508, new_AGEMA_signal_19505, new_AGEMA_signal_19502}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_8138, new_AGEMA_signal_8137, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_19517, new_AGEMA_signal_19514, new_AGEMA_signal_19511}), .clk (clk), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_8120, new_AGEMA_signal_8119, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_19526, new_AGEMA_signal_19523, new_AGEMA_signal_19520}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_19535, new_AGEMA_signal_19532, new_AGEMA_signal_19529}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_19544, new_AGEMA_signal_19541, new_AGEMA_signal_19538}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_8126, new_AGEMA_signal_8125, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_8138, new_AGEMA_signal_8137, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_8132, new_AGEMA_signal_8131, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9830, new_AGEMA_signal_9829, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9836, new_AGEMA_signal_9835, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9842, new_AGEMA_signal_9841, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9836, new_AGEMA_signal_9835, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_9830, new_AGEMA_signal_9829, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_9842, new_AGEMA_signal_9841, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_19553, new_AGEMA_signal_19550, new_AGEMA_signal_19547}), .clk (clk), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_19562, new_AGEMA_signal_19559, new_AGEMA_signal_19556}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_8150, new_AGEMA_signal_8149, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_19571, new_AGEMA_signal_19568, new_AGEMA_signal_19565}), .clk (clk), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_19580, new_AGEMA_signal_19577, new_AGEMA_signal_19574}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_19589, new_AGEMA_signal_19586, new_AGEMA_signal_19583}), .clk (clk), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_19598, new_AGEMA_signal_19595, new_AGEMA_signal_19592}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_19607, new_AGEMA_signal_19604, new_AGEMA_signal_19601}), .clk (clk), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_19616, new_AGEMA_signal_19613, new_AGEMA_signal_19610}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_19625, new_AGEMA_signal_19622, new_AGEMA_signal_19619}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_19634, new_AGEMA_signal_19631, new_AGEMA_signal_19628}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_19643, new_AGEMA_signal_19640, new_AGEMA_signal_19637}), .clk (clk), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_19652, new_AGEMA_signal_19649, new_AGEMA_signal_19646}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_19661, new_AGEMA_signal_19658, new_AGEMA_signal_19655}), .clk (clk), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_19670, new_AGEMA_signal_19667, new_AGEMA_signal_19664}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_19679, new_AGEMA_signal_19676, new_AGEMA_signal_19673}), .clk (clk), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_8144, new_AGEMA_signal_8143, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_19688, new_AGEMA_signal_19685, new_AGEMA_signal_19682}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_19697, new_AGEMA_signal_19694, new_AGEMA_signal_19691}), .clk (clk), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_19706, new_AGEMA_signal_19703, new_AGEMA_signal_19700}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_8150, new_AGEMA_signal_8149, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_8156, new_AGEMA_signal_8155, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9854, new_AGEMA_signal_9853, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9482, new_AGEMA_signal_9481, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9860, new_AGEMA_signal_9859, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_8642, new_AGEMA_signal_8641, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_9854, new_AGEMA_signal_9853, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_9860, new_AGEMA_signal_9859, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9482, new_AGEMA_signal_9481, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_19715, new_AGEMA_signal_19712, new_AGEMA_signal_19709}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_19724, new_AGEMA_signal_19721, new_AGEMA_signal_19718}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_19733, new_AGEMA_signal_19730, new_AGEMA_signal_19727}), .clk (clk), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_19742, new_AGEMA_signal_19739, new_AGEMA_signal_19736}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_19751, new_AGEMA_signal_19748, new_AGEMA_signal_19745}), .clk (clk), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_19760, new_AGEMA_signal_19757, new_AGEMA_signal_19754}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_19769, new_AGEMA_signal_19766, new_AGEMA_signal_19763}), .clk (clk), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_19778, new_AGEMA_signal_19775, new_AGEMA_signal_19772}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_19787, new_AGEMA_signal_19784, new_AGEMA_signal_19781}), .clk (clk), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_8654, new_AGEMA_signal_8653, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_19796, new_AGEMA_signal_19793, new_AGEMA_signal_19790}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_19805, new_AGEMA_signal_19802, new_AGEMA_signal_19799}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_19814, new_AGEMA_signal_19811, new_AGEMA_signal_19808}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_19823, new_AGEMA_signal_19820, new_AGEMA_signal_19817}), .clk (clk), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_19832, new_AGEMA_signal_19829, new_AGEMA_signal_19826}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_19841, new_AGEMA_signal_19838, new_AGEMA_signal_19835}), .clk (clk), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_19850, new_AGEMA_signal_19847, new_AGEMA_signal_19844}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_19859, new_AGEMA_signal_19856, new_AGEMA_signal_19853}), .clk (clk), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_19868, new_AGEMA_signal_19865, new_AGEMA_signal_19862}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_8654, new_AGEMA_signal_8653, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_8648, new_AGEMA_signal_8647, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_8660, new_AGEMA_signal_8659, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9500, new_AGEMA_signal_9499, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_9488, new_AGEMA_signal_9487, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_8666, new_AGEMA_signal_8665, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_9494, new_AGEMA_signal_9493, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9500, new_AGEMA_signal_9499, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_19877, new_AGEMA_signal_19874, new_AGEMA_signal_19871}), .clk (clk), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_19886, new_AGEMA_signal_19883, new_AGEMA_signal_19880}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_19895, new_AGEMA_signal_19892, new_AGEMA_signal_19889}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_19904, new_AGEMA_signal_19901, new_AGEMA_signal_19898}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_19913, new_AGEMA_signal_19910, new_AGEMA_signal_19907}), .clk (clk), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_19922, new_AGEMA_signal_19919, new_AGEMA_signal_19916}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_19931, new_AGEMA_signal_19928, new_AGEMA_signal_19925}), .clk (clk), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_19940, new_AGEMA_signal_19937, new_AGEMA_signal_19934}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_19949, new_AGEMA_signal_19946, new_AGEMA_signal_19943}), .clk (clk), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_8678, new_AGEMA_signal_8677, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_19958, new_AGEMA_signal_19955, new_AGEMA_signal_19952}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_19967, new_AGEMA_signal_19964, new_AGEMA_signal_19961}), .clk (clk), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_19976, new_AGEMA_signal_19973, new_AGEMA_signal_19970}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_19985, new_AGEMA_signal_19982, new_AGEMA_signal_19979}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_19994, new_AGEMA_signal_19991, new_AGEMA_signal_19988}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_20003, new_AGEMA_signal_20000, new_AGEMA_signal_19997}), .clk (clk), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_20012, new_AGEMA_signal_20009, new_AGEMA_signal_20006}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_20021, new_AGEMA_signal_20018, new_AGEMA_signal_20015}), .clk (clk), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_20030, new_AGEMA_signal_20027, new_AGEMA_signal_20024}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_8678, new_AGEMA_signal_8677, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_8672, new_AGEMA_signal_8671, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_8684, new_AGEMA_signal_8683, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_9518, new_AGEMA_signal_9517, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_9506, new_AGEMA_signal_9505, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_9512, new_AGEMA_signal_9511, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_9518, new_AGEMA_signal_9517, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_20039, new_AGEMA_signal_20036, new_AGEMA_signal_20033}), .clk (clk), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_20048, new_AGEMA_signal_20045, new_AGEMA_signal_20042}), .clk (clk), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_20057, new_AGEMA_signal_20054, new_AGEMA_signal_20051}), .clk (clk), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_20066, new_AGEMA_signal_20063, new_AGEMA_signal_20060}), .clk (clk), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_20075, new_AGEMA_signal_20072, new_AGEMA_signal_20069}), .clk (clk), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_20084, new_AGEMA_signal_20081, new_AGEMA_signal_20078}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_20093, new_AGEMA_signal_20090, new_AGEMA_signal_20087}), .clk (clk), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_20102, new_AGEMA_signal_20099, new_AGEMA_signal_20096}), .clk (clk), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_20111, new_AGEMA_signal_20108, new_AGEMA_signal_20105}), .clk (clk), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_20120, new_AGEMA_signal_20117, new_AGEMA_signal_20114}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_20129, new_AGEMA_signal_20126, new_AGEMA_signal_20123}), .clk (clk), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_20138, new_AGEMA_signal_20135, new_AGEMA_signal_20132}), .clk (clk), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_20147, new_AGEMA_signal_20144, new_AGEMA_signal_20141}), .clk (clk), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_20156, new_AGEMA_signal_20153, new_AGEMA_signal_20150}), .clk (clk), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_20165, new_AGEMA_signal_20162, new_AGEMA_signal_20159}), .clk (clk), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_20174, new_AGEMA_signal_20171, new_AGEMA_signal_20168}), .clk (clk), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_20183, new_AGEMA_signal_20180, new_AGEMA_signal_20177}), .clk (clk), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_20192, new_AGEMA_signal_20189, new_AGEMA_signal_20186}), .clk (clk), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_9524, new_AGEMA_signal_9523, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_20201, new_AGEMA_signal_20198, new_AGEMA_signal_20195}), .clk (clk), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_20210, new_AGEMA_signal_20207, new_AGEMA_signal_20204}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_20219, new_AGEMA_signal_20216, new_AGEMA_signal_20213}), .clk (clk), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_20228, new_AGEMA_signal_20225, new_AGEMA_signal_20222}), .clk (clk), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_20237, new_AGEMA_signal_20234, new_AGEMA_signal_20231}), .clk (clk), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_20246, new_AGEMA_signal_20243, new_AGEMA_signal_20240}), .clk (clk), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_20255, new_AGEMA_signal_20252, new_AGEMA_signal_20249}), .clk (clk), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_20264, new_AGEMA_signal_20261, new_AGEMA_signal_20258}), .clk (clk), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_20273, new_AGEMA_signal_20270, new_AGEMA_signal_20267}), .clk (clk), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_20282, new_AGEMA_signal_20279, new_AGEMA_signal_20276}), .clk (clk), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_20291, new_AGEMA_signal_20288, new_AGEMA_signal_20285}), .clk (clk), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_20300, new_AGEMA_signal_20297, new_AGEMA_signal_20294}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_20309, new_AGEMA_signal_20306, new_AGEMA_signal_20303}), .clk (clk), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_20318, new_AGEMA_signal_20315, new_AGEMA_signal_20312}), .clk (clk), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_20327, new_AGEMA_signal_20324, new_AGEMA_signal_20321}), .clk (clk), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_20336, new_AGEMA_signal_20333, new_AGEMA_signal_20330}), .clk (clk), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_20345, new_AGEMA_signal_20342, new_AGEMA_signal_20339}), .clk (clk), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_20354, new_AGEMA_signal_20351, new_AGEMA_signal_20348}), .clk (clk), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_20363, new_AGEMA_signal_20360, new_AGEMA_signal_20357}), .clk (clk), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_20372, new_AGEMA_signal_20369, new_AGEMA_signal_20366}), .clk (clk), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_20381, new_AGEMA_signal_20378, new_AGEMA_signal_20375}), .clk (clk), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_20390, new_AGEMA_signal_20387, new_AGEMA_signal_20384}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_20399, new_AGEMA_signal_20396, new_AGEMA_signal_20393}), .clk (clk), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_20408, new_AGEMA_signal_20405, new_AGEMA_signal_20402}), .clk (clk), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_20417, new_AGEMA_signal_20414, new_AGEMA_signal_20411}), .clk (clk), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_20426, new_AGEMA_signal_20423, new_AGEMA_signal_20420}), .clk (clk), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_20435, new_AGEMA_signal_20432, new_AGEMA_signal_20429}), .clk (clk), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_20444, new_AGEMA_signal_20441, new_AGEMA_signal_20438}), .clk (clk), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_20453, new_AGEMA_signal_20450, new_AGEMA_signal_20447}), .clk (clk), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_20462, new_AGEMA_signal_20459, new_AGEMA_signal_20456}), .clk (clk), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_20471, new_AGEMA_signal_20468, new_AGEMA_signal_20465}), .clk (clk), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_20480, new_AGEMA_signal_20477, new_AGEMA_signal_20474}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_20489, new_AGEMA_signal_20486, new_AGEMA_signal_20483}), .clk (clk), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_20498, new_AGEMA_signal_20495, new_AGEMA_signal_20492}), .clk (clk), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_20507, new_AGEMA_signal_20504, new_AGEMA_signal_20501}), .clk (clk), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_20516, new_AGEMA_signal_20513, new_AGEMA_signal_20510}), .clk (clk), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_9188, new_AGEMA_signal_9187, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_9188, new_AGEMA_signal_9187, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9194, new_AGEMA_signal_9193, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_9182, new_AGEMA_signal_9181, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_9194, new_AGEMA_signal_9193, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_20525, new_AGEMA_signal_20522, new_AGEMA_signal_20519}), .clk (clk), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_20534, new_AGEMA_signal_20531, new_AGEMA_signal_20528}), .clk (clk), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_20543, new_AGEMA_signal_20540, new_AGEMA_signal_20537}), .clk (clk), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_20552, new_AGEMA_signal_20549, new_AGEMA_signal_20546}), .clk (clk), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_20561, new_AGEMA_signal_20558, new_AGEMA_signal_20555}), .clk (clk), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_20570, new_AGEMA_signal_20567, new_AGEMA_signal_20564}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_20579, new_AGEMA_signal_20576, new_AGEMA_signal_20573}), .clk (clk), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_20588, new_AGEMA_signal_20585, new_AGEMA_signal_20582}), .clk (clk), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_20597, new_AGEMA_signal_20594, new_AGEMA_signal_20591}), .clk (clk), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_20606, new_AGEMA_signal_20603, new_AGEMA_signal_20600}), .clk (clk), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_20615, new_AGEMA_signal_20612, new_AGEMA_signal_20609}), .clk (clk), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_20624, new_AGEMA_signal_20621, new_AGEMA_signal_20618}), .clk (clk), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_20633, new_AGEMA_signal_20630, new_AGEMA_signal_20627}), .clk (clk), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_20642, new_AGEMA_signal_20639, new_AGEMA_signal_20636}), .clk (clk), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_20651, new_AGEMA_signal_20648, new_AGEMA_signal_20645}), .clk (clk), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_20660, new_AGEMA_signal_20657, new_AGEMA_signal_20654}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_20669, new_AGEMA_signal_20666, new_AGEMA_signal_20663}), .clk (clk), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_20678, new_AGEMA_signal_20675, new_AGEMA_signal_20672}), .clk (clk), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_9200, new_AGEMA_signal_9199, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9212, new_AGEMA_signal_9211, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_9206, new_AGEMA_signal_9205, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_9212, new_AGEMA_signal_9211, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_20687, new_AGEMA_signal_20684, new_AGEMA_signal_20681}), .clk (clk), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_20696, new_AGEMA_signal_20693, new_AGEMA_signal_20690}), .clk (clk), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_20705, new_AGEMA_signal_20702, new_AGEMA_signal_20699}), .clk (clk), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_20714, new_AGEMA_signal_20711, new_AGEMA_signal_20708}), .clk (clk), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_20723, new_AGEMA_signal_20720, new_AGEMA_signal_20717}), .clk (clk), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_20732, new_AGEMA_signal_20729, new_AGEMA_signal_20726}), .clk (clk), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_20741, new_AGEMA_signal_20738, new_AGEMA_signal_20735}), .clk (clk), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_20750, new_AGEMA_signal_20747, new_AGEMA_signal_20744}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_20759, new_AGEMA_signal_20756, new_AGEMA_signal_20753}), .clk (clk), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_20768, new_AGEMA_signal_20765, new_AGEMA_signal_20762}), .clk (clk), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_20777, new_AGEMA_signal_20774, new_AGEMA_signal_20771}), .clk (clk), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_20786, new_AGEMA_signal_20783, new_AGEMA_signal_20780}), .clk (clk), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_20795, new_AGEMA_signal_20792, new_AGEMA_signal_20789}), .clk (clk), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_20804, new_AGEMA_signal_20801, new_AGEMA_signal_20798}), .clk (clk), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_20813, new_AGEMA_signal_20810, new_AGEMA_signal_20807}), .clk (clk), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_20822, new_AGEMA_signal_20819, new_AGEMA_signal_20816}), .clk (clk), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_20831, new_AGEMA_signal_20828, new_AGEMA_signal_20825}), .clk (clk), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_20840, new_AGEMA_signal_20837, new_AGEMA_signal_20834}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_9218, new_AGEMA_signal_9217, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_9230, new_AGEMA_signal_9229, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_9236, new_AGEMA_signal_9235, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_9224, new_AGEMA_signal_9223, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_9236, new_AGEMA_signal_9235, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_9230, new_AGEMA_signal_9229, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_20849, new_AGEMA_signal_20846, new_AGEMA_signal_20843}), .clk (clk), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_20858, new_AGEMA_signal_20855, new_AGEMA_signal_20852}), .clk (clk), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_20867, new_AGEMA_signal_20864, new_AGEMA_signal_20861}), .clk (clk), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_20876, new_AGEMA_signal_20873, new_AGEMA_signal_20870}), .clk (clk), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_20885, new_AGEMA_signal_20882, new_AGEMA_signal_20879}), .clk (clk), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_20894, new_AGEMA_signal_20891, new_AGEMA_signal_20888}), .clk (clk), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_20903, new_AGEMA_signal_20900, new_AGEMA_signal_20897}), .clk (clk), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_20912, new_AGEMA_signal_20909, new_AGEMA_signal_20906}), .clk (clk), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_20921, new_AGEMA_signal_20918, new_AGEMA_signal_20915}), .clk (clk), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_20930, new_AGEMA_signal_20927, new_AGEMA_signal_20924}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_20939, new_AGEMA_signal_20936, new_AGEMA_signal_20933}), .clk (clk), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_20948, new_AGEMA_signal_20945, new_AGEMA_signal_20942}), .clk (clk), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_20957, new_AGEMA_signal_20954, new_AGEMA_signal_20951}), .clk (clk), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_20966, new_AGEMA_signal_20963, new_AGEMA_signal_20960}), .clk (clk), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_20975, new_AGEMA_signal_20972, new_AGEMA_signal_20969}), .clk (clk), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_20984, new_AGEMA_signal_20981, new_AGEMA_signal_20978}), .clk (clk), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_20993, new_AGEMA_signal_20990, new_AGEMA_signal_20987}), .clk (clk), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_21002, new_AGEMA_signal_20999, new_AGEMA_signal_20996}), .clk (clk), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_21011, new_AGEMA_signal_21008, new_AGEMA_signal_21005}), .clk (clk), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_21020, new_AGEMA_signal_21017, new_AGEMA_signal_21014}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_21029, new_AGEMA_signal_21026, new_AGEMA_signal_21023}), .clk (clk), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_21038, new_AGEMA_signal_21035, new_AGEMA_signal_21032}), .clk (clk), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_21047, new_AGEMA_signal_21044, new_AGEMA_signal_21041}), .clk (clk), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_21056, new_AGEMA_signal_21053, new_AGEMA_signal_21050}), .clk (clk), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_21065, new_AGEMA_signal_21062, new_AGEMA_signal_21059}), .clk (clk), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_21074, new_AGEMA_signal_21071, new_AGEMA_signal_21068}), .clk (clk), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_21083, new_AGEMA_signal_21080, new_AGEMA_signal_21077}), .clk (clk), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_21092, new_AGEMA_signal_21089, new_AGEMA_signal_21086}), .clk (clk), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_21101, new_AGEMA_signal_21098, new_AGEMA_signal_21095}), .clk (clk), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_21110, new_AGEMA_signal_21107, new_AGEMA_signal_21104}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_21119, new_AGEMA_signal_21116, new_AGEMA_signal_21113}), .clk (clk), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_21128, new_AGEMA_signal_21125, new_AGEMA_signal_21122}), .clk (clk), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_21137, new_AGEMA_signal_21134, new_AGEMA_signal_21131}), .clk (clk), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_21146, new_AGEMA_signal_21143, new_AGEMA_signal_21140}), .clk (clk), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_21155, new_AGEMA_signal_21152, new_AGEMA_signal_21149}), .clk (clk), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_21164, new_AGEMA_signal_21161, new_AGEMA_signal_21158}), .clk (clk), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_21173, new_AGEMA_signal_21170, new_AGEMA_signal_21167}), .clk (clk), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_21182, new_AGEMA_signal_21179, new_AGEMA_signal_21176}), .clk (clk), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_21191, new_AGEMA_signal_21188, new_AGEMA_signal_21185}), .clk (clk), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_21200, new_AGEMA_signal_21197, new_AGEMA_signal_21194}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_21209, new_AGEMA_signal_21206, new_AGEMA_signal_21203}), .clk (clk), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_21218, new_AGEMA_signal_21215, new_AGEMA_signal_21212}), .clk (clk), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_21227, new_AGEMA_signal_21224, new_AGEMA_signal_21221}), .clk (clk), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_21236, new_AGEMA_signal_21233, new_AGEMA_signal_21230}), .clk (clk), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_21245, new_AGEMA_signal_21242, new_AGEMA_signal_21239}), .clk (clk), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_21254, new_AGEMA_signal_21251, new_AGEMA_signal_21248}), .clk (clk), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_21263, new_AGEMA_signal_21260, new_AGEMA_signal_21257}), .clk (clk), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_21272, new_AGEMA_signal_21269, new_AGEMA_signal_21266}), .clk (clk), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_21281, new_AGEMA_signal_21278, new_AGEMA_signal_21275}), .clk (clk), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_21290, new_AGEMA_signal_21287, new_AGEMA_signal_21284}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({new_AGEMA_signal_8402, new_AGEMA_signal_8401, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_21299, new_AGEMA_signal_21296, new_AGEMA_signal_21293}), .clk (clk), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_21308, new_AGEMA_signal_21305, new_AGEMA_signal_21302}), .clk (clk), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_21317, new_AGEMA_signal_21314, new_AGEMA_signal_21311}), .clk (clk), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_21326, new_AGEMA_signal_21323, new_AGEMA_signal_21320}), .clk (clk), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_8402, new_AGEMA_signal_8401, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_8882, new_AGEMA_signal_8881, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_21335, new_AGEMA_signal_21332, new_AGEMA_signal_21329}), .clk (clk), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_21344, new_AGEMA_signal_21341, new_AGEMA_signal_21338}), .clk (clk), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({new_AGEMA_signal_8414, new_AGEMA_signal_8413, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_21353, new_AGEMA_signal_21350, new_AGEMA_signal_21347}), .clk (clk), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_21362, new_AGEMA_signal_21359, new_AGEMA_signal_21356}), .clk (clk), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_21371, new_AGEMA_signal_21368, new_AGEMA_signal_21365}), .clk (clk), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_21380, new_AGEMA_signal_21377, new_AGEMA_signal_21374}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_21389, new_AGEMA_signal_21386, new_AGEMA_signal_21383}), .clk (clk), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_21398, new_AGEMA_signal_21395, new_AGEMA_signal_21392}), .clk (clk), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_21407, new_AGEMA_signal_21404, new_AGEMA_signal_21401}), .clk (clk), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_8894, new_AGEMA_signal_8893, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_21416, new_AGEMA_signal_21413, new_AGEMA_signal_21410}), .clk (clk), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_21425, new_AGEMA_signal_21422, new_AGEMA_signal_21419}), .clk (clk), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_21434, new_AGEMA_signal_21431, new_AGEMA_signal_21428}), .clk (clk), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_21443, new_AGEMA_signal_21440, new_AGEMA_signal_21437}), .clk (clk), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_21452, new_AGEMA_signal_21449, new_AGEMA_signal_21446}), .clk (clk), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({new_AGEMA_signal_8426, new_AGEMA_signal_8425, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_21461, new_AGEMA_signal_21458, new_AGEMA_signal_21455}), .clk (clk), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_8408, new_AGEMA_signal_8407, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_21470, new_AGEMA_signal_21467, new_AGEMA_signal_21464}), .clk (clk), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_21479, new_AGEMA_signal_21476, new_AGEMA_signal_21473}), .clk (clk), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_21488, new_AGEMA_signal_21485, new_AGEMA_signal_21482}), .clk (clk), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_8414, new_AGEMA_signal_8413, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_8894, new_AGEMA_signal_8893, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_8888, new_AGEMA_signal_8887, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_8426, new_AGEMA_signal_8425, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_8420, new_AGEMA_signal_8419, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_8900, new_AGEMA_signal_8899, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_8906, new_AGEMA_signal_8905, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_21497, new_AGEMA_signal_21494, new_AGEMA_signal_21491}), .clk (clk), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_21506, new_AGEMA_signal_21503, new_AGEMA_signal_21500}), .clk (clk), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({new_AGEMA_signal_8438, new_AGEMA_signal_8437, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_21515, new_AGEMA_signal_21512, new_AGEMA_signal_21509}), .clk (clk), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_21524, new_AGEMA_signal_21521, new_AGEMA_signal_21518}), .clk (clk), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_21533, new_AGEMA_signal_21530, new_AGEMA_signal_21527}), .clk (clk), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_21542, new_AGEMA_signal_21539, new_AGEMA_signal_21536}), .clk (clk), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_21551, new_AGEMA_signal_21548, new_AGEMA_signal_21545}), .clk (clk), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_21560, new_AGEMA_signal_21557, new_AGEMA_signal_21554}), .clk (clk), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_21569, new_AGEMA_signal_21566, new_AGEMA_signal_21563}), .clk (clk), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({new_AGEMA_signal_8918, new_AGEMA_signal_8917, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_21578, new_AGEMA_signal_21575, new_AGEMA_signal_21572}), .clk (clk), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_21587, new_AGEMA_signal_21584, new_AGEMA_signal_21581}), .clk (clk), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_21596, new_AGEMA_signal_21593, new_AGEMA_signal_21590}), .clk (clk), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_21605, new_AGEMA_signal_21602, new_AGEMA_signal_21599}), .clk (clk), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_21614, new_AGEMA_signal_21611, new_AGEMA_signal_21608}), .clk (clk), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_21623, new_AGEMA_signal_21620, new_AGEMA_signal_21617}), .clk (clk), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_8432, new_AGEMA_signal_8431, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_21632, new_AGEMA_signal_21629, new_AGEMA_signal_21626}), .clk (clk), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_21641, new_AGEMA_signal_21638, new_AGEMA_signal_21635}), .clk (clk), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_21650, new_AGEMA_signal_21647, new_AGEMA_signal_21644}), .clk (clk), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_8438, new_AGEMA_signal_8437, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_8918, new_AGEMA_signal_8917, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_8912, new_AGEMA_signal_8911, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_8444, new_AGEMA_signal_8443, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_8924, new_AGEMA_signal_8923, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_8930, new_AGEMA_signal_8929, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_21659, new_AGEMA_signal_21656, new_AGEMA_signal_21653}), .clk (clk), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_21668, new_AGEMA_signal_21665, new_AGEMA_signal_21662}), .clk (clk), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_21677, new_AGEMA_signal_21674, new_AGEMA_signal_21671}), .clk (clk), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_21686, new_AGEMA_signal_21683, new_AGEMA_signal_21680}), .clk (clk), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_21695, new_AGEMA_signal_21692, new_AGEMA_signal_21689}), .clk (clk), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_21704, new_AGEMA_signal_21701, new_AGEMA_signal_21698}), .clk (clk), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_21713, new_AGEMA_signal_21710, new_AGEMA_signal_21707}), .clk (clk), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_21722, new_AGEMA_signal_21719, new_AGEMA_signal_21716}), .clk (clk), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_21731, new_AGEMA_signal_21728, new_AGEMA_signal_21725}), .clk (clk), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_21740, new_AGEMA_signal_21737, new_AGEMA_signal_21734}), .clk (clk), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_21749, new_AGEMA_signal_21746, new_AGEMA_signal_21743}), .clk (clk), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_21758, new_AGEMA_signal_21755, new_AGEMA_signal_21752}), .clk (clk), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_21767, new_AGEMA_signal_21764, new_AGEMA_signal_21761}), .clk (clk), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_21776, new_AGEMA_signal_21773, new_AGEMA_signal_21770}), .clk (clk), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_21785, new_AGEMA_signal_21782, new_AGEMA_signal_21779}), .clk (clk), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_21794, new_AGEMA_signal_21791, new_AGEMA_signal_21788}), .clk (clk), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_21803, new_AGEMA_signal_21800, new_AGEMA_signal_21797}), .clk (clk), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_21812, new_AGEMA_signal_21809, new_AGEMA_signal_21806}), .clk (clk), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_8936, new_AGEMA_signal_8935, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_11390, new_AGEMA_signal_11389, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, MixColumnsOutput[105]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_11390, new_AGEMA_signal_11389, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, MixColumnsOutput[104]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .c ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, MixColumnsOutput[103]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_10946, new_AGEMA_signal_10945, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_11396, new_AGEMA_signal_11395, MixColumnsOutput[102]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_10946, new_AGEMA_signal_10945, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, MixColumnsOutput[101]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, MixColumnsOutput[100]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_11402, new_AGEMA_signal_11401, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_11996, new_AGEMA_signal_11995, MixColumnsOutput[99]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .c ({new_AGEMA_signal_11402, new_AGEMA_signal_11401, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, MixColumnsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_10952, new_AGEMA_signal_10951, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, MixColumnsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_10952, new_AGEMA_signal_10951, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_11408, new_AGEMA_signal_11407, MixColumnsOutput[98]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .c ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, MixColumnsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_10526, new_AGEMA_signal_10525, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, MixColumnsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_10562, new_AGEMA_signal_10561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_10958, new_AGEMA_signal_10957, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_11414, new_AGEMA_signal_11413, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, MixColumnsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .b ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .b ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_11414, new_AGEMA_signal_11413, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, MixColumnsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_12002, new_AGEMA_signal_12001, MixColumnsOutput[121]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_10964, new_AGEMA_signal_10963, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_11420, new_AGEMA_signal_11419, MixColumnsOutput[120]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10964, new_AGEMA_signal_10963, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, MixColumnsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, MixColumnsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_10532, new_AGEMA_signal_10531, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_10970, new_AGEMA_signal_10969, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_11426, new_AGEMA_signal_11425, MixColumnsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_10970, new_AGEMA_signal_10969, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, MixColumnsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_10568, new_AGEMA_signal_10567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, MixColumnsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_10976, new_AGEMA_signal_10975, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_11432, new_AGEMA_signal_11431, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_12008, new_AGEMA_signal_12007, MixColumnsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .b ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_11432, new_AGEMA_signal_11431, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, MixColumnsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .b ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .b ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, MixColumnsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_10982, new_AGEMA_signal_10981, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_11438, new_AGEMA_signal_11437, MixColumnsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_10538, new_AGEMA_signal_10537, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_10988, new_AGEMA_signal_10987, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, MixColumnsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_10988, new_AGEMA_signal_10987, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_10544, new_AGEMA_signal_10543, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, MixColumnsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_10364, new_AGEMA_signal_10363, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_11444, new_AGEMA_signal_11443, MixColumnsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_10226, new_AGEMA_signal_10225, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_10298, new_AGEMA_signal_10297, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_10550, new_AGEMA_signal_10549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10436, new_AGEMA_signal_10435, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, MixColumnsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_10574, new_AGEMA_signal_10573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_10994, new_AGEMA_signal_10993, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_10580, new_AGEMA_signal_10579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_12014, new_AGEMA_signal_12013, MixColumnsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .b ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .c ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .c ({new_AGEMA_signal_11000, new_AGEMA_signal_10999, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_11450, new_AGEMA_signal_11449, MixColumnsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .b ({new_AGEMA_signal_10304, new_AGEMA_signal_10303, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .c ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .c ({new_AGEMA_signal_10556, new_AGEMA_signal_10555, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .c ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, MixColumnsOutput[96]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .c ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, MixColumnsInput[123]}), .c ({new_AGEMA_signal_10562, new_AGEMA_signal_10561, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10442, new_AGEMA_signal_10441, MixColumnsInput[122]}), .c ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, MixColumnsInput[120]}), .c ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10370, new_AGEMA_signal_10369, MixColumnsInput[115]}), .c ({new_AGEMA_signal_10568, new_AGEMA_signal_10567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, MixColumnsInput[114]}), .c ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_10046, new_AGEMA_signal_10045, MixColumnsInput[112]}), .c ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, MixColumnsInput[107]}), .c ({new_AGEMA_signal_10574, new_AGEMA_signal_10573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, MixColumnsInput[106]}), .c ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10292, new_AGEMA_signal_10291, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, MixColumnsInput[104]}), .c ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, MixColumnsInput[99]}), .c ({new_AGEMA_signal_10580, new_AGEMA_signal_10579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_10232, new_AGEMA_signal_10231, MixColumnsInput[98]}), .c ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, MixColumnsInput[96]}), .c ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, MixColumnsOutput[73]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_11006, new_AGEMA_signal_11005, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_11456, new_AGEMA_signal_11455, MixColumnsOutput[72]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .c ({new_AGEMA_signal_11006, new_AGEMA_signal_11005, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, MixColumnsOutput[71]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, MixColumnsOutput[70]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_11012, new_AGEMA_signal_11011, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_11462, new_AGEMA_signal_11461, MixColumnsOutput[69]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_11012, new_AGEMA_signal_11011, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, MixColumnsOutput[68]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_12020, new_AGEMA_signal_12019, MixColumnsOutput[67]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .c ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_11468, new_AGEMA_signal_11467, MixColumnsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_10586, new_AGEMA_signal_10585, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, MixColumnsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_11018, new_AGEMA_signal_11017, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, MixColumnsOutput[66]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .c ({new_AGEMA_signal_11018, new_AGEMA_signal_11017, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_11474, new_AGEMA_signal_11473, MixColumnsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, MixColumnsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, MixColumnsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .b ({new_AGEMA_signal_10628, new_AGEMA_signal_10627, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_11024, new_AGEMA_signal_11023, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .b ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_11480, new_AGEMA_signal_11479, MixColumnsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_10592, new_AGEMA_signal_10591, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .b ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_12026, new_AGEMA_signal_12025, MixColumnsOutput[89]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, MixColumnsOutput[88]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_11030, new_AGEMA_signal_11029, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_11486, new_AGEMA_signal_11485, MixColumnsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_11030, new_AGEMA_signal_11029, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, MixColumnsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, MixColumnsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_10598, new_AGEMA_signal_10597, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_11492, new_AGEMA_signal_11491, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, MixColumnsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_11036, new_AGEMA_signal_11035, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_11492, new_AGEMA_signal_11491, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, MixColumnsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_12032, new_AGEMA_signal_12031, MixColumnsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .b ({new_AGEMA_signal_10634, new_AGEMA_signal_10633, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_11042, new_AGEMA_signal_11041, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .b ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_11498, new_AGEMA_signal_11497, MixColumnsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .b ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, MixColumnsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_10388, new_AGEMA_signal_10387, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_11048, new_AGEMA_signal_11047, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, MixColumnsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .b ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_10604, new_AGEMA_signal_10603, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_11504, new_AGEMA_signal_11503, MixColumnsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10238, new_AGEMA_signal_10237, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_11054, new_AGEMA_signal_11053, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, MixColumnsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_10610, new_AGEMA_signal_10609, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_11054, new_AGEMA_signal_11053, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, MixColumnsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_10394, new_AGEMA_signal_10393, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_10310, new_AGEMA_signal_10309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_10616, new_AGEMA_signal_10615, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_11510, new_AGEMA_signal_11509, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, MixColumnsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_11510, new_AGEMA_signal_11509, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_10382, new_AGEMA_signal_10381, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_11060, new_AGEMA_signal_11059, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_12038, new_AGEMA_signal_12037, MixColumnsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .b ({new_AGEMA_signal_10640, new_AGEMA_signal_10639, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .c ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_10646, new_AGEMA_signal_10645, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .c ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_11066, new_AGEMA_signal_11065, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, MixColumnsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .c ({new_AGEMA_signal_11066, new_AGEMA_signal_11065, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .c ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .c ({new_AGEMA_signal_11516, new_AGEMA_signal_11515, MixColumnsOutput[64]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .b ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_10622, new_AGEMA_signal_10621, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .c ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, MixColumnsInput[91]}), .c ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, MixColumnsInput[90]}), .c ({new_AGEMA_signal_10628, new_AGEMA_signal_10627, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10376, new_AGEMA_signal_10375, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, MixColumnsInput[88]}), .c ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, MixColumnsInput[83]}), .c ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_10316, new_AGEMA_signal_10315, MixColumnsInput[82]}), .c ({new_AGEMA_signal_10634, new_AGEMA_signal_10633, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, MixColumnsInput[80]}), .c ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10244, new_AGEMA_signal_10243, MixColumnsInput[75]}), .c ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, MixColumnsInput[74]}), .c ({new_AGEMA_signal_10640, new_AGEMA_signal_10639, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_9848, new_AGEMA_signal_9847, MixColumnsInput[72]}), .c ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, MixColumnsInput[67]}), .c ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10400, new_AGEMA_signal_10399, MixColumnsInput[66]}), .c ({new_AGEMA_signal_10646, new_AGEMA_signal_10645, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, MixColumnsInput[64]}), .c ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, MixColumnsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, MixColumnsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .c ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_11072, new_AGEMA_signal_11071, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_11522, new_AGEMA_signal_11521, MixColumnsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_11072, new_AGEMA_signal_11071, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, MixColumnsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, MixColumnsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_11528, new_AGEMA_signal_11527, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, MixColumnsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_11528, new_AGEMA_signal_11527, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_12044, new_AGEMA_signal_12043, MixColumnsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .c ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_11078, new_AGEMA_signal_11077, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, MixColumnsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_11078, new_AGEMA_signal_11077, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_11534, new_AGEMA_signal_11533, MixColumnsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_10652, new_AGEMA_signal_10651, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, MixColumnsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .c ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_11084, new_AGEMA_signal_11083, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, MixColumnsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_11084, new_AGEMA_signal_11083, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_11540, new_AGEMA_signal_11539, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, MixColumnsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_11540, new_AGEMA_signal_11539, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, MixColumnsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .b ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_11090, new_AGEMA_signal_11089, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, MixColumnsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .b ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_11090, new_AGEMA_signal_11089, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_11546, new_AGEMA_signal_11545, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_12050, new_AGEMA_signal_12049, MixColumnsOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_11546, new_AGEMA_signal_11545, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, MixColumnsOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, MixColumnsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_10658, new_AGEMA_signal_10657, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_11096, new_AGEMA_signal_11095, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_11552, new_AGEMA_signal_11551, MixColumnsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_11096, new_AGEMA_signal_11095, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, MixColumnsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, MixColumnsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_11558, new_AGEMA_signal_11557, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, MixColumnsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_10694, new_AGEMA_signal_10693, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_11102, new_AGEMA_signal_11101, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_11558, new_AGEMA_signal_11557, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_10712, new_AGEMA_signal_10711, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_12056, new_AGEMA_signal_12055, MixColumnsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .b ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .b ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_11108, new_AGEMA_signal_11107, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, MixColumnsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .b ({new_AGEMA_signal_10262, new_AGEMA_signal_10261, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_10664, new_AGEMA_signal_10663, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .b ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_11108, new_AGEMA_signal_11107, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_11564, new_AGEMA_signal_11563, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, MixColumnsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_10700, new_AGEMA_signal_10699, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_11564, new_AGEMA_signal_11563, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_10706, new_AGEMA_signal_10705, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_11114, new_AGEMA_signal_11113, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, MixColumnsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .b ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_11114, new_AGEMA_signal_11113, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, MixColumnsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10406, new_AGEMA_signal_10405, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_10670, new_AGEMA_signal_10669, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_11570, new_AGEMA_signal_11569, MixColumnsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10322, new_AGEMA_signal_10321, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_10676, new_AGEMA_signal_10675, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_11120, new_AGEMA_signal_11119, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, MixColumnsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_11120, new_AGEMA_signal_11119, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, MixColumnsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_10340, new_AGEMA_signal_10339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_10256, new_AGEMA_signal_10255, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_11576, new_AGEMA_signal_11575, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_12062, new_AGEMA_signal_12061, MixColumnsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .b ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_11126, new_AGEMA_signal_11125, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .c ({new_AGEMA_signal_11576, new_AGEMA_signal_11575, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .c ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, MixColumnsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .b ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_10682, new_AGEMA_signal_10681, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .c ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_10346, new_AGEMA_signal_10345, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .c ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_11132, new_AGEMA_signal_11131, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .c ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, MixColumnsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_11132, new_AGEMA_signal_11131, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .c ({new_AGEMA_signal_10688, new_AGEMA_signal_10687, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10328, new_AGEMA_signal_10327, MixColumnsInput[59]}), .c ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, MixColumnsInput[58]}), .c ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_9980, new_AGEMA_signal_9979, MixColumnsInput[56]}), .c ({new_AGEMA_signal_10694, new_AGEMA_signal_10693, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, MixColumnsInput[51]}), .c ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, MixColumnsInput[50]}), .c ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10250, new_AGEMA_signal_10249, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, MixColumnsInput[48]}), .c ({new_AGEMA_signal_10700, new_AGEMA_signal_10699, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10412, new_AGEMA_signal_10411, MixColumnsInput[43]}), .c ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, MixColumnsInput[42]}), .c ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_10112, new_AGEMA_signal_10111, MixColumnsInput[40]}), .c ({new_AGEMA_signal_10706, new_AGEMA_signal_10705, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, MixColumnsInput[35]}), .c ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, MixColumnsInput[34]}), .c ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10334, new_AGEMA_signal_10333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, MixColumnsInput[32]}), .c ({new_AGEMA_signal_10712, new_AGEMA_signal_10711, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_11582, new_AGEMA_signal_11581, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_11582, new_AGEMA_signal_11581, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .c ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_11138, new_AGEMA_signal_11137, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_11588, new_AGEMA_signal_11587, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_11138, new_AGEMA_signal_11137, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_11594, new_AGEMA_signal_11593, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_12068, new_AGEMA_signal_12067, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .c ({new_AGEMA_signal_11594, new_AGEMA_signal_11593, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_11144, new_AGEMA_signal_11143, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_11144, new_AGEMA_signal_11143, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_11600, new_AGEMA_signal_11599, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .c ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_10718, new_AGEMA_signal_10717, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_10754, new_AGEMA_signal_10753, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_11150, new_AGEMA_signal_11149, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_11606, new_AGEMA_signal_11605, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .b ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .b ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_11606, new_AGEMA_signal_11605, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_12074, new_AGEMA_signal_12073, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_11156, new_AGEMA_signal_11155, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_11612, new_AGEMA_signal_11611, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_11156, new_AGEMA_signal_11155, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_10724, new_AGEMA_signal_10723, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_11162, new_AGEMA_signal_11161, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_11618, new_AGEMA_signal_11617, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_11162, new_AGEMA_signal_11161, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_10760, new_AGEMA_signal_10759, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_11168, new_AGEMA_signal_11167, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_11624, new_AGEMA_signal_11623, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_12080, new_AGEMA_signal_12079, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .b ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .b ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_11624, new_AGEMA_signal_11623, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .b ({new_AGEMA_signal_10430, new_AGEMA_signal_10429, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_11174, new_AGEMA_signal_11173, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_11630, new_AGEMA_signal_11629, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_10730, new_AGEMA_signal_10729, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .b ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_11180, new_AGEMA_signal_11179, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_11180, new_AGEMA_signal_11179, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_10736, new_AGEMA_signal_10735, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_10280, new_AGEMA_signal_10279, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_10352, new_AGEMA_signal_10351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_11636, new_AGEMA_signal_11635, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_10742, new_AGEMA_signal_10741, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_10268, new_AGEMA_signal_10267, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_10766, new_AGEMA_signal_10765, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_11186, new_AGEMA_signal_11185, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_10424, new_AGEMA_signal_10423, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_10772, new_AGEMA_signal_10771, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_12086, new_AGEMA_signal_12085, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .b ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .c ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .c ({new_AGEMA_signal_11192, new_AGEMA_signal_11191, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_11642, new_AGEMA_signal_11641, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .b ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .c ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .c ({new_AGEMA_signal_10748, new_AGEMA_signal_10747, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .c ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .c ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, MixColumnsInput[27]}), .c ({new_AGEMA_signal_10754, new_AGEMA_signal_10753, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_10274, new_AGEMA_signal_10273, MixColumnsInput[26]}), .c ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, MixColumnsInput[24]}), .c ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, MixColumnsInput[19]}), .c ({new_AGEMA_signal_10760, new_AGEMA_signal_10759, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, MixColumnsInput[18]}), .c ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_10418, new_AGEMA_signal_10417, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, MixColumnsInput[16]}), .c ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, MixColumnsInput[11]}), .c ({new_AGEMA_signal_10766, new_AGEMA_signal_10765, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10358, new_AGEMA_signal_10357, MixColumnsInput[10]}), .c ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, MixColumnsInput[8]}), .c ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10286, new_AGEMA_signal_10285, MixColumnsInput[3]}), .c ({new_AGEMA_signal_10772, new_AGEMA_signal_10771, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, MixColumnsInput[2]}), .c ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_9914, new_AGEMA_signal_9913, MixColumnsInput[0]}), .c ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, KeyExpansionOutput[0]}), .a ({new_AGEMA_signal_21824, new_AGEMA_signal_21820, new_AGEMA_signal_21816}), .c ({new_AGEMA_signal_11648, new_AGEMA_signal_11647, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, KeyExpansionOutput[1]}), .a ({new_AGEMA_signal_21836, new_AGEMA_signal_21832, new_AGEMA_signal_21828}), .c ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, KeyExpansionOutput[2]}), .a ({new_AGEMA_signal_21848, new_AGEMA_signal_21844, new_AGEMA_signal_21840}), .c ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, KeyExpansionOutput[3]}), .a ({new_AGEMA_signal_21860, new_AGEMA_signal_21856, new_AGEMA_signal_21852}), .c ({new_AGEMA_signal_12098, new_AGEMA_signal_12097, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, KeyExpansionOutput[4]}), .a ({new_AGEMA_signal_21872, new_AGEMA_signal_21868, new_AGEMA_signal_21864}), .c ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionOutput[5]}), .a ({new_AGEMA_signal_21884, new_AGEMA_signal_21880, new_AGEMA_signal_21876}), .c ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, KeyExpansionOutput[6]}), .a ({new_AGEMA_signal_21896, new_AGEMA_signal_21892, new_AGEMA_signal_21888}), .c ({new_AGEMA_signal_12110, new_AGEMA_signal_12109, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, KeyExpansionOutput[7]}), .a ({new_AGEMA_signal_21908, new_AGEMA_signal_21904, new_AGEMA_signal_21900}), .c ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, KeyExpansionOutput[8]}), .a ({new_AGEMA_signal_21920, new_AGEMA_signal_21916, new_AGEMA_signal_21912}), .c ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionOutput[9]}), .a ({new_AGEMA_signal_21932, new_AGEMA_signal_21928, new_AGEMA_signal_21924}), .c ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, KeyExpansionOutput[10]}), .a ({new_AGEMA_signal_21944, new_AGEMA_signal_21940, new_AGEMA_signal_21936}), .c ({new_AGEMA_signal_12122, new_AGEMA_signal_12121, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionOutput[11]}), .a ({new_AGEMA_signal_21956, new_AGEMA_signal_21952, new_AGEMA_signal_21948}), .c ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, KeyExpansionOutput[12]}), .a ({new_AGEMA_signal_21968, new_AGEMA_signal_21964, new_AGEMA_signal_21960}), .c ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, KeyExpansionOutput[13]}), .a ({new_AGEMA_signal_21980, new_AGEMA_signal_21976, new_AGEMA_signal_21972}), .c ({new_AGEMA_signal_12134, new_AGEMA_signal_12133, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionOutput[14]}), .a ({new_AGEMA_signal_21992, new_AGEMA_signal_21988, new_AGEMA_signal_21984}), .c ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, KeyExpansionOutput[15]}), .a ({new_AGEMA_signal_22004, new_AGEMA_signal_22000, new_AGEMA_signal_21996}), .c ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, KeyExpansionOutput[16]}), .a ({new_AGEMA_signal_22016, new_AGEMA_signal_22012, new_AGEMA_signal_22008}), .c ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, KeyExpansionOutput[17]}), .a ({new_AGEMA_signal_22028, new_AGEMA_signal_22024, new_AGEMA_signal_22020}), .c ({new_AGEMA_signal_12146, new_AGEMA_signal_12145, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionOutput[18]}), .a ({new_AGEMA_signal_22040, new_AGEMA_signal_22036, new_AGEMA_signal_22032}), .c ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, KeyExpansionOutput[19]}), .a ({new_AGEMA_signal_22052, new_AGEMA_signal_22048, new_AGEMA_signal_22044}), .c ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionOutput[20]}), .a ({new_AGEMA_signal_22064, new_AGEMA_signal_22060, new_AGEMA_signal_22056}), .c ({new_AGEMA_signal_12158, new_AGEMA_signal_12157, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, KeyExpansionOutput[21]}), .a ({new_AGEMA_signal_22076, new_AGEMA_signal_22072, new_AGEMA_signal_22068}), .c ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, KeyExpansionOutput[22]}), .a ({new_AGEMA_signal_22088, new_AGEMA_signal_22084, new_AGEMA_signal_22080}), .c ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionOutput[23]}), .a ({new_AGEMA_signal_22100, new_AGEMA_signal_22096, new_AGEMA_signal_22092}), .c ({new_AGEMA_signal_12170, new_AGEMA_signal_12169, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, KeyExpansionOutput[24]}), .a ({new_AGEMA_signal_22112, new_AGEMA_signal_22108, new_AGEMA_signal_22104}), .c ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, KeyExpansionOutput[25]}), .a ({new_AGEMA_signal_22124, new_AGEMA_signal_22120, new_AGEMA_signal_22116}), .c ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, KeyExpansionOutput[26]}), .a ({new_AGEMA_signal_22136, new_AGEMA_signal_22132, new_AGEMA_signal_22128}), .c ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12212, new_AGEMA_signal_12211, KeyExpansionOutput[27]}), .a ({new_AGEMA_signal_22148, new_AGEMA_signal_22144, new_AGEMA_signal_22140}), .c ({new_AGEMA_signal_12644, new_AGEMA_signal_12643, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, KeyExpansionOutput[28]}), .a ({new_AGEMA_signal_22160, new_AGEMA_signal_22156, new_AGEMA_signal_22152}), .c ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, KeyExpansionOutput[29]}), .a ({new_AGEMA_signal_22172, new_AGEMA_signal_22168, new_AGEMA_signal_22164}), .c ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12206, new_AGEMA_signal_12205, KeyExpansionOutput[30]}), .a ({new_AGEMA_signal_22184, new_AGEMA_signal_22180, new_AGEMA_signal_22176}), .c ({new_AGEMA_signal_12656, new_AGEMA_signal_12655, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, KeyExpansionOutput[31]}), .a ({new_AGEMA_signal_22196, new_AGEMA_signal_22192, new_AGEMA_signal_22188}), .c ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}), .a ({new_AGEMA_signal_22208, new_AGEMA_signal_22204, new_AGEMA_signal_22200}), .c ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}), .a ({new_AGEMA_signal_22220, new_AGEMA_signal_22216, new_AGEMA_signal_22212}), .c ({new_AGEMA_signal_11660, new_AGEMA_signal_11659, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}), .a ({new_AGEMA_signal_22232, new_AGEMA_signal_22228, new_AGEMA_signal_22224}), .c ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}), .a ({new_AGEMA_signal_22244, new_AGEMA_signal_22240, new_AGEMA_signal_22236}), .c ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}), .a ({new_AGEMA_signal_22256, new_AGEMA_signal_22252, new_AGEMA_signal_22248}), .c ({new_AGEMA_signal_11672, new_AGEMA_signal_11671, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}), .a ({new_AGEMA_signal_22268, new_AGEMA_signal_22264, new_AGEMA_signal_22260}), .c ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}), .a ({new_AGEMA_signal_22280, new_AGEMA_signal_22276, new_AGEMA_signal_22272}), .c ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}), .a ({new_AGEMA_signal_22292, new_AGEMA_signal_22288, new_AGEMA_signal_22284}), .c ({new_AGEMA_signal_11684, new_AGEMA_signal_11683, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}), .a ({new_AGEMA_signal_22304, new_AGEMA_signal_22300, new_AGEMA_signal_22296}), .c ({new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}), .a ({new_AGEMA_signal_22316, new_AGEMA_signal_22312, new_AGEMA_signal_22308}), .c ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}), .a ({new_AGEMA_signal_22328, new_AGEMA_signal_22324, new_AGEMA_signal_22320}), .c ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}), .a ({new_AGEMA_signal_22340, new_AGEMA_signal_22336, new_AGEMA_signal_22332}), .c ({new_AGEMA_signal_11696, new_AGEMA_signal_11695, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}), .a ({new_AGEMA_signal_22352, new_AGEMA_signal_22348, new_AGEMA_signal_22344}), .c ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}), .a ({new_AGEMA_signal_22364, new_AGEMA_signal_22360, new_AGEMA_signal_22356}), .c ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}), .a ({new_AGEMA_signal_22376, new_AGEMA_signal_22372, new_AGEMA_signal_22368}), .c ({new_AGEMA_signal_11708, new_AGEMA_signal_11707, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}), .a ({new_AGEMA_signal_22388, new_AGEMA_signal_22384, new_AGEMA_signal_22380}), .c ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}), .a ({new_AGEMA_signal_22400, new_AGEMA_signal_22396, new_AGEMA_signal_22392}), .c ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}), .a ({new_AGEMA_signal_22412, new_AGEMA_signal_22408, new_AGEMA_signal_22404}), .c ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}), .a ({new_AGEMA_signal_22424, new_AGEMA_signal_22420, new_AGEMA_signal_22416}), .c ({new_AGEMA_signal_11720, new_AGEMA_signal_11719, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}), .a ({new_AGEMA_signal_22436, new_AGEMA_signal_22432, new_AGEMA_signal_22428}), .c ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}), .a ({new_AGEMA_signal_22448, new_AGEMA_signal_22444, new_AGEMA_signal_22440}), .c ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}), .a ({new_AGEMA_signal_22460, new_AGEMA_signal_22456, new_AGEMA_signal_22452}), .c ({new_AGEMA_signal_11732, new_AGEMA_signal_11731, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}), .a ({new_AGEMA_signal_22472, new_AGEMA_signal_22468, new_AGEMA_signal_22464}), .c ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}), .a ({new_AGEMA_signal_22484, new_AGEMA_signal_22480, new_AGEMA_signal_22476}), .c ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}), .a ({new_AGEMA_signal_22496, new_AGEMA_signal_22492, new_AGEMA_signal_22488}), .c ({new_AGEMA_signal_11744, new_AGEMA_signal_11743, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}), .a ({new_AGEMA_signal_22508, new_AGEMA_signal_22504, new_AGEMA_signal_22500}), .c ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}), .a ({new_AGEMA_signal_22520, new_AGEMA_signal_22516, new_AGEMA_signal_22512}), .c ({new_AGEMA_signal_12182, new_AGEMA_signal_12181, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}), .a ({new_AGEMA_signal_22532, new_AGEMA_signal_22528, new_AGEMA_signal_22524}), .c ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}), .a ({new_AGEMA_signal_22544, new_AGEMA_signal_22540, new_AGEMA_signal_22536}), .c ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}), .a ({new_AGEMA_signal_22556, new_AGEMA_signal_22552, new_AGEMA_signal_22548}), .c ({new_AGEMA_signal_12194, new_AGEMA_signal_12193, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}), .a ({new_AGEMA_signal_22568, new_AGEMA_signal_22564, new_AGEMA_signal_22560}), .c ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}), .a ({new_AGEMA_signal_22580, new_AGEMA_signal_22576, new_AGEMA_signal_22572}), .c ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}), .a ({new_AGEMA_signal_22592, new_AGEMA_signal_22588, new_AGEMA_signal_22584}), .c ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}), .a ({new_AGEMA_signal_22604, new_AGEMA_signal_22600, new_AGEMA_signal_22596}), .c ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}), .a ({new_AGEMA_signal_22616, new_AGEMA_signal_22612, new_AGEMA_signal_22608}), .c ({new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}), .a ({new_AGEMA_signal_22628, new_AGEMA_signal_22624, new_AGEMA_signal_22620}), .c ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}), .a ({new_AGEMA_signal_22640, new_AGEMA_signal_22636, new_AGEMA_signal_22632}), .c ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}), .a ({new_AGEMA_signal_22652, new_AGEMA_signal_22648, new_AGEMA_signal_22644}), .c ({new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}), .a ({new_AGEMA_signal_22664, new_AGEMA_signal_22660, new_AGEMA_signal_22656}), .c ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}), .a ({new_AGEMA_signal_22676, new_AGEMA_signal_22672, new_AGEMA_signal_22668}), .c ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}), .a ({new_AGEMA_signal_22688, new_AGEMA_signal_22684, new_AGEMA_signal_22680}), .c ({new_AGEMA_signal_10784, new_AGEMA_signal_10783, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}), .a ({new_AGEMA_signal_22700, new_AGEMA_signal_22696, new_AGEMA_signal_22692}), .c ({new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}), .a ({new_AGEMA_signal_22712, new_AGEMA_signal_22708, new_AGEMA_signal_22704}), .c ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}), .a ({new_AGEMA_signal_22724, new_AGEMA_signal_22720, new_AGEMA_signal_22716}), .c ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}), .a ({new_AGEMA_signal_22736, new_AGEMA_signal_22732, new_AGEMA_signal_22728}), .c ({new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}), .a ({new_AGEMA_signal_22748, new_AGEMA_signal_22744, new_AGEMA_signal_22740}), .c ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}), .a ({new_AGEMA_signal_22760, new_AGEMA_signal_22756, new_AGEMA_signal_22752}), .c ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}), .a ({new_AGEMA_signal_22772, new_AGEMA_signal_22768, new_AGEMA_signal_22764}), .c ({new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}), .a ({new_AGEMA_signal_22784, new_AGEMA_signal_22780, new_AGEMA_signal_22776}), .c ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}), .a ({new_AGEMA_signal_22796, new_AGEMA_signal_22792, new_AGEMA_signal_22788}), .c ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}), .a ({new_AGEMA_signal_22808, new_AGEMA_signal_22804, new_AGEMA_signal_22800}), .c ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}), .a ({new_AGEMA_signal_22820, new_AGEMA_signal_22816, new_AGEMA_signal_22812}), .c ({new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}), .a ({new_AGEMA_signal_22832, new_AGEMA_signal_22828, new_AGEMA_signal_22824}), .c ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}), .a ({new_AGEMA_signal_22844, new_AGEMA_signal_22840, new_AGEMA_signal_22836}), .c ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}), .a ({new_AGEMA_signal_22856, new_AGEMA_signal_22852, new_AGEMA_signal_22848}), .c ({new_AGEMA_signal_11288, new_AGEMA_signal_11287, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}), .a ({new_AGEMA_signal_22868, new_AGEMA_signal_22864, new_AGEMA_signal_22860}), .c ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}), .a ({new_AGEMA_signal_22880, new_AGEMA_signal_22876, new_AGEMA_signal_22872}), .c ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}), .a ({new_AGEMA_signal_22892, new_AGEMA_signal_22888, new_AGEMA_signal_22884}), .c ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}), .a ({new_AGEMA_signal_22904, new_AGEMA_signal_22900, new_AGEMA_signal_22896}), .c ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}), .a ({new_AGEMA_signal_22916, new_AGEMA_signal_22912, new_AGEMA_signal_22908}), .c ({new_AGEMA_signal_11756, new_AGEMA_signal_11755, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}), .a ({new_AGEMA_signal_22928, new_AGEMA_signal_22924, new_AGEMA_signal_22920}), .c ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}), .a ({new_AGEMA_signal_22940, new_AGEMA_signal_22936, new_AGEMA_signal_22932}), .c ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}), .a ({new_AGEMA_signal_22952, new_AGEMA_signal_22948, new_AGEMA_signal_22944}), .c ({new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}), .a ({new_AGEMA_signal_22964, new_AGEMA_signal_22960, new_AGEMA_signal_22956}), .c ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}), .a ({new_AGEMA_signal_22976, new_AGEMA_signal_22972, new_AGEMA_signal_22968}), .c ({new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}), .a ({new_AGEMA_signal_22988, new_AGEMA_signal_22984, new_AGEMA_signal_22980}), .c ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}), .a ({new_AGEMA_signal_23000, new_AGEMA_signal_22996, new_AGEMA_signal_22992}), .c ({new_AGEMA_signal_10796, new_AGEMA_signal_10795, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}), .a ({new_AGEMA_signal_23012, new_AGEMA_signal_23008, new_AGEMA_signal_23004}), .c ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}), .a ({new_AGEMA_signal_23024, new_AGEMA_signal_23020, new_AGEMA_signal_23016}), .c ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}), .a ({new_AGEMA_signal_23036, new_AGEMA_signal_23032, new_AGEMA_signal_23028}), .c ({new_AGEMA_signal_10808, new_AGEMA_signal_10807, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}), .a ({new_AGEMA_signal_23048, new_AGEMA_signal_23044, new_AGEMA_signal_23040}), .c ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}), .a ({new_AGEMA_signal_23060, new_AGEMA_signal_23056, new_AGEMA_signal_23052}), .c ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}), .a ({new_AGEMA_signal_23072, new_AGEMA_signal_23068, new_AGEMA_signal_23064}), .c ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}), .a ({new_AGEMA_signal_23084, new_AGEMA_signal_23080, new_AGEMA_signal_23076}), .c ({new_AGEMA_signal_10820, new_AGEMA_signal_10819, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}), .a ({new_AGEMA_signal_23096, new_AGEMA_signal_23092, new_AGEMA_signal_23088}), .c ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}), .a ({new_AGEMA_signal_23108, new_AGEMA_signal_23104, new_AGEMA_signal_23100}), .c ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}), .a ({new_AGEMA_signal_23120, new_AGEMA_signal_23116, new_AGEMA_signal_23112}), .c ({new_AGEMA_signal_10832, new_AGEMA_signal_10831, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}), .a ({new_AGEMA_signal_23132, new_AGEMA_signal_23128, new_AGEMA_signal_23124}), .c ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}), .a ({new_AGEMA_signal_23144, new_AGEMA_signal_23140, new_AGEMA_signal_23136}), .c ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}), .a ({new_AGEMA_signal_23156, new_AGEMA_signal_23152, new_AGEMA_signal_23148}), .c ({new_AGEMA_signal_10844, new_AGEMA_signal_10843, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}), .a ({new_AGEMA_signal_23168, new_AGEMA_signal_23164, new_AGEMA_signal_23160}), .c ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}), .a ({new_AGEMA_signal_23180, new_AGEMA_signal_23176, new_AGEMA_signal_23172}), .c ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}), .a ({new_AGEMA_signal_23192, new_AGEMA_signal_23188, new_AGEMA_signal_23184}), .c ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}), .a ({new_AGEMA_signal_23204, new_AGEMA_signal_23200, new_AGEMA_signal_23196}), .c ({new_AGEMA_signal_10856, new_AGEMA_signal_10855, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}), .a ({new_AGEMA_signal_23216, new_AGEMA_signal_23212, new_AGEMA_signal_23208}), .c ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}), .a ({new_AGEMA_signal_23228, new_AGEMA_signal_23224, new_AGEMA_signal_23220}), .c ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}), .a ({new_AGEMA_signal_23240, new_AGEMA_signal_23236, new_AGEMA_signal_23232}), .c ({new_AGEMA_signal_10868, new_AGEMA_signal_10867, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}), .a ({new_AGEMA_signal_23252, new_AGEMA_signal_23248, new_AGEMA_signal_23244}), .c ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}), .a ({new_AGEMA_signal_23264, new_AGEMA_signal_23260, new_AGEMA_signal_23256}), .c ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}), .a ({new_AGEMA_signal_23276, new_AGEMA_signal_23272, new_AGEMA_signal_23268}), .c ({new_AGEMA_signal_11300, new_AGEMA_signal_11299, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}), .a ({new_AGEMA_signal_23288, new_AGEMA_signal_23284, new_AGEMA_signal_23280}), .c ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}), .a ({new_AGEMA_signal_23300, new_AGEMA_signal_23296, new_AGEMA_signal_23292}), .c ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}), .a ({new_AGEMA_signal_23312, new_AGEMA_signal_23308, new_AGEMA_signal_23304}), .c ({new_AGEMA_signal_11312, new_AGEMA_signal_11311, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}), .a ({new_AGEMA_signal_23324, new_AGEMA_signal_23320, new_AGEMA_signal_23316}), .c ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}), .a ({new_AGEMA_signal_23336, new_AGEMA_signal_23332, new_AGEMA_signal_23328}), .c ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_17684), .b ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}), .a ({new_AGEMA_signal_23348, new_AGEMA_signal_23344, new_AGEMA_signal_23340}), .c ({new_AGEMA_signal_11324, new_AGEMA_signal_11323, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_23360, new_AGEMA_signal_23356, new_AGEMA_signal_23352}), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_23372, new_AGEMA_signal_23368, new_AGEMA_signal_23364}), .b ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_23384, new_AGEMA_signal_23380, new_AGEMA_signal_23376}), .b ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_23396, new_AGEMA_signal_23392, new_AGEMA_signal_23388}), .b ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_23408, new_AGEMA_signal_23404, new_AGEMA_signal_23400}), .b ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_23420, new_AGEMA_signal_23416, new_AGEMA_signal_23412}), .b ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_23432, new_AGEMA_signal_23428, new_AGEMA_signal_23424}), .b ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_23444, new_AGEMA_signal_23440, new_AGEMA_signal_23436}), .b ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_23456, new_AGEMA_signal_23452, new_AGEMA_signal_23448}), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_10880, new_AGEMA_signal_10879, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_23468, new_AGEMA_signal_23464, new_AGEMA_signal_23460}), .b ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_23480, new_AGEMA_signal_23476, new_AGEMA_signal_23472}), .b ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_23492, new_AGEMA_signal_23488, new_AGEMA_signal_23484}), .b ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_11330, new_AGEMA_signal_11329, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_23504, new_AGEMA_signal_23500, new_AGEMA_signal_23496}), .b ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_23516, new_AGEMA_signal_23512, new_AGEMA_signal_23508}), .b ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_23528, new_AGEMA_signal_23524, new_AGEMA_signal_23520}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_23540, new_AGEMA_signal_23536, new_AGEMA_signal_23532}), .b ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_23552, new_AGEMA_signal_23548, new_AGEMA_signal_23544}), .b ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_10886, new_AGEMA_signal_10885, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_23564, new_AGEMA_signal_23560, new_AGEMA_signal_23556}), .b ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_11336, new_AGEMA_signal_11335, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_23576, new_AGEMA_signal_23572, new_AGEMA_signal_23568}), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_23588, new_AGEMA_signal_23584, new_AGEMA_signal_23580}), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_23600, new_AGEMA_signal_23596, new_AGEMA_signal_23592}), .b ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_23612, new_AGEMA_signal_23608, new_AGEMA_signal_23604}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_23624, new_AGEMA_signal_23620, new_AGEMA_signal_23616}), .b ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_23636, new_AGEMA_signal_23632, new_AGEMA_signal_23628}), .b ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_23648, new_AGEMA_signal_23644, new_AGEMA_signal_23640}), .b ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_23660, new_AGEMA_signal_23656, new_AGEMA_signal_23652}), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_12206, new_AGEMA_signal_12205, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_23672, new_AGEMA_signal_23668, new_AGEMA_signal_23664}), .b ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_23684, new_AGEMA_signal_23680, new_AGEMA_signal_23676}), .b ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_11342, new_AGEMA_signal_11341, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_23696, new_AGEMA_signal_23692, new_AGEMA_signal_23688}), .b ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_23708, new_AGEMA_signal_23704, new_AGEMA_signal_23700}), .b ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_23720, new_AGEMA_signal_23716, new_AGEMA_signal_23712}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_10892, new_AGEMA_signal_10891, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_23732, new_AGEMA_signal_23728, new_AGEMA_signal_23724}), .b ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_23744, new_AGEMA_signal_23740, new_AGEMA_signal_23736}), .b ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_23756, new_AGEMA_signal_23752, new_AGEMA_signal_23748}), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_23768, new_AGEMA_signal_23764, new_AGEMA_signal_23760}), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_23780, new_AGEMA_signal_23776, new_AGEMA_signal_23772}), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_23792, new_AGEMA_signal_23788, new_AGEMA_signal_23784}), .b ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_23804, new_AGEMA_signal_23800, new_AGEMA_signal_23796}), .b ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_11348, new_AGEMA_signal_11347, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_23816, new_AGEMA_signal_23812, new_AGEMA_signal_23808}), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_12212, new_AGEMA_signal_12211, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_23828, new_AGEMA_signal_23824, new_AGEMA_signal_23820}), .b ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_23840, new_AGEMA_signal_23836, new_AGEMA_signal_23832}), .b ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_23852, new_AGEMA_signal_23848, new_AGEMA_signal_23844}), .b ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_23864, new_AGEMA_signal_23860, new_AGEMA_signal_23856}), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_23876, new_AGEMA_signal_23872, new_AGEMA_signal_23868}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_23888, new_AGEMA_signal_23884, new_AGEMA_signal_23880}), .b ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_23900, new_AGEMA_signal_23896, new_AGEMA_signal_23892}), .b ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_23912, new_AGEMA_signal_23908, new_AGEMA_signal_23904}), .b ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_11354, new_AGEMA_signal_11353, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_23924, new_AGEMA_signal_23920, new_AGEMA_signal_23916}), .b ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_23936, new_AGEMA_signal_23932, new_AGEMA_signal_23928}), .b ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_23948, new_AGEMA_signal_23944, new_AGEMA_signal_23940}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_23960, new_AGEMA_signal_23956, new_AGEMA_signal_23952}), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_23972, new_AGEMA_signal_23968, new_AGEMA_signal_23964}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_23984, new_AGEMA_signal_23980, new_AGEMA_signal_23976}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_23996, new_AGEMA_signal_23992, new_AGEMA_signal_23988}), .b ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_24008, new_AGEMA_signal_24004, new_AGEMA_signal_24000}), .b ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_11360, new_AGEMA_signal_11359, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_24020, new_AGEMA_signal_24016, new_AGEMA_signal_24012}), .b ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_10898, new_AGEMA_signal_10897, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_24032, new_AGEMA_signal_24028, new_AGEMA_signal_24024}), .b ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_24044, new_AGEMA_signal_24040, new_AGEMA_signal_24036}), .b ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_24056, new_AGEMA_signal_24052, new_AGEMA_signal_24048}), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_24068, new_AGEMA_signal_24064, new_AGEMA_signal_24060}), .b ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_24080, new_AGEMA_signal_24076, new_AGEMA_signal_24072}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_24092, new_AGEMA_signal_24088, new_AGEMA_signal_24084}), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_24104, new_AGEMA_signal_24100, new_AGEMA_signal_24096}), .b ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_24116, new_AGEMA_signal_24112, new_AGEMA_signal_24108}), .b ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_11366, new_AGEMA_signal_11365, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_24128, new_AGEMA_signal_24124, new_AGEMA_signal_24120}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_10904, new_AGEMA_signal_10903, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_24140, new_AGEMA_signal_24136, new_AGEMA_signal_24132}), .b ({new_AGEMA_signal_10220, new_AGEMA_signal_10219, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_24152, new_AGEMA_signal_24148, new_AGEMA_signal_24144}), .b ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_24164, new_AGEMA_signal_24160, new_AGEMA_signal_24156}), .b ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_24176, new_AGEMA_signal_24172, new_AGEMA_signal_24168}), .b ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_24188, new_AGEMA_signal_24184, new_AGEMA_signal_24180}), .b ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_24200, new_AGEMA_signal_24196, new_AGEMA_signal_24192}), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_24212, new_AGEMA_signal_24208, new_AGEMA_signal_24204}), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_24224, new_AGEMA_signal_24220, new_AGEMA_signal_24216}), .b ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_24236, new_AGEMA_signal_24232, new_AGEMA_signal_24228}), .b ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_11372, new_AGEMA_signal_11371, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_24248, new_AGEMA_signal_24244, new_AGEMA_signal_24240}), .b ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_10910, new_AGEMA_signal_10909, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_24260, new_AGEMA_signal_24256, new_AGEMA_signal_24252}), .b ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_24272, new_AGEMA_signal_24268, new_AGEMA_signal_24264}), .b ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_24284, new_AGEMA_signal_24280, new_AGEMA_signal_24276}), .b ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_24296, new_AGEMA_signal_24292, new_AGEMA_signal_24288}), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_24308, new_AGEMA_signal_24304, new_AGEMA_signal_24300}), .b ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_24320, new_AGEMA_signal_24316, new_AGEMA_signal_24312}), .b ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_24332, new_AGEMA_signal_24328, new_AGEMA_signal_24324}), .b ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_24344, new_AGEMA_signal_24340, new_AGEMA_signal_24336}), .b ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_11378, new_AGEMA_signal_11377, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_24356, new_AGEMA_signal_24352, new_AGEMA_signal_24348}), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_10916, new_AGEMA_signal_10915, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_24368, new_AGEMA_signal_24364, new_AGEMA_signal_24360}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_24380, new_AGEMA_signal_24376, new_AGEMA_signal_24372}), .b ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_24392, new_AGEMA_signal_24388, new_AGEMA_signal_24384}), .b ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_24404, new_AGEMA_signal_24400, new_AGEMA_signal_24396}), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_24416, new_AGEMA_signal_24412, new_AGEMA_signal_24408}), .b ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_24428, new_AGEMA_signal_24424, new_AGEMA_signal_24420}), .b ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_24440, new_AGEMA_signal_24436, new_AGEMA_signal_24432}), .b ({new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_10922, new_AGEMA_signal_10921, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_24452, new_AGEMA_signal_24448, new_AGEMA_signal_24444}), .b ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_24464, new_AGEMA_signal_24460, new_AGEMA_signal_24456}), .b ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_24476, new_AGEMA_signal_24472, new_AGEMA_signal_24468}), .b ({new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_10928, new_AGEMA_signal_10927, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_24488, new_AGEMA_signal_24484, new_AGEMA_signal_24480}), .b ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_24500, new_AGEMA_signal_24496, new_AGEMA_signal_24492}), .b ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_24512, new_AGEMA_signal_24508, new_AGEMA_signal_24504}), .b ({new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_10934, new_AGEMA_signal_10933, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_24524, new_AGEMA_signal_24520, new_AGEMA_signal_24516}), .b ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_24536, new_AGEMA_signal_24532, new_AGEMA_signal_24528}), .b ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_24548, new_AGEMA_signal_24544, new_AGEMA_signal_24540}), .b ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_11384, new_AGEMA_signal_11383, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_24560, new_AGEMA_signal_24556, new_AGEMA_signal_24552}), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_24572, new_AGEMA_signal_24568, new_AGEMA_signal_24564}), .b ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_24584, new_AGEMA_signal_24580, new_AGEMA_signal_24576}), .b ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_24596, new_AGEMA_signal_24592, new_AGEMA_signal_24588}), .b ({new_AGEMA_signal_10184, new_AGEMA_signal_10183, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_24608, new_AGEMA_signal_24604, new_AGEMA_signal_24600}), .b ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_24620, new_AGEMA_signal_24616, new_AGEMA_signal_24612}), .b ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_24632, new_AGEMA_signal_24628, new_AGEMA_signal_24624}), .b ({new_AGEMA_signal_10190, new_AGEMA_signal_10189, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_24644, new_AGEMA_signal_24640, new_AGEMA_signal_24636}), .b ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_24656, new_AGEMA_signal_24652, new_AGEMA_signal_24648}), .b ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_24668, new_AGEMA_signal_24664, new_AGEMA_signal_24660}), .b ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_24680, new_AGEMA_signal_24676, new_AGEMA_signal_24672}), .b ({new_AGEMA_signal_10196, new_AGEMA_signal_10195, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_24692, new_AGEMA_signal_24688, new_AGEMA_signal_24684}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_24704, new_AGEMA_signal_24700, new_AGEMA_signal_24696}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_24716, new_AGEMA_signal_24712, new_AGEMA_signal_24708}), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_24728, new_AGEMA_signal_24724, new_AGEMA_signal_24720}), .b ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_24740, new_AGEMA_signal_24736, new_AGEMA_signal_24732}), .b ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_24752, new_AGEMA_signal_24748, new_AGEMA_signal_24744}), .b ({new_AGEMA_signal_10202, new_AGEMA_signal_10201, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_24764, new_AGEMA_signal_24760, new_AGEMA_signal_24756}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_24776, new_AGEMA_signal_24772, new_AGEMA_signal_24768}), .b ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_24788, new_AGEMA_signal_24784, new_AGEMA_signal_24780}), .b ({new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_10160, new_AGEMA_signal_10159, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_24800, new_AGEMA_signal_24796, new_AGEMA_signal_24792}), .b ({new_AGEMA_signal_10208, new_AGEMA_signal_10207, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_24812, new_AGEMA_signal_24808, new_AGEMA_signal_24804}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_24824, new_AGEMA_signal_24820, new_AGEMA_signal_24816}), .b ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_24836, new_AGEMA_signal_24832, new_AGEMA_signal_24828}), .b ({new_AGEMA_signal_10214, new_AGEMA_signal_10213, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_24848, new_AGEMA_signal_24844, new_AGEMA_signal_24840}), .b ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_24860, new_AGEMA_signal_24856, new_AGEMA_signal_24852}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_10940, new_AGEMA_signal_10939, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_24872, new_AGEMA_signal_24868, new_AGEMA_signal_24864}), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_24884, new_AGEMA_signal_24880, new_AGEMA_signal_24876}), .b ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_10166, new_AGEMA_signal_10165, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24888}), .c ({new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24892}), .c ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24896}), .c ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_10172, new_AGEMA_signal_10171, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24900}), .c ({new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24904}), .c ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24908}), .c ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_10178, new_AGEMA_signal_10177, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24912}), .c ({new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, 1'b0, new_AGEMA_signal_24916}), .c ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_24925, new_AGEMA_signal_24922, new_AGEMA_signal_24919}), .clk (clk), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_24934, new_AGEMA_signal_24931, new_AGEMA_signal_24928}), .clk (clk), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({new_AGEMA_signal_8006, new_AGEMA_signal_8005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_24259, new_AGEMA_signal_24255, new_AGEMA_signal_24251}), .clk (clk), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_24943, new_AGEMA_signal_24940, new_AGEMA_signal_24937}), .clk (clk), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_24952, new_AGEMA_signal_24949, new_AGEMA_signal_24946}), .clk (clk), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_24961, new_AGEMA_signal_24958, new_AGEMA_signal_24955}), .clk (clk), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_24970, new_AGEMA_signal_24967, new_AGEMA_signal_24964}), .clk (clk), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_24979, new_AGEMA_signal_24976, new_AGEMA_signal_24973}), .clk (clk), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_24988, new_AGEMA_signal_24985, new_AGEMA_signal_24982}), .clk (clk), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({new_AGEMA_signal_8486, new_AGEMA_signal_8485, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_24997, new_AGEMA_signal_24994, new_AGEMA_signal_24991}), .clk (clk), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_7844, new_AGEMA_signal_7843, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_25006, new_AGEMA_signal_25003, new_AGEMA_signal_25000}), .clk (clk), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_25015, new_AGEMA_signal_25012, new_AGEMA_signal_25009}), .clk (clk), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_25024, new_AGEMA_signal_25021, new_AGEMA_signal_25018}), .clk (clk), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_25033, new_AGEMA_signal_25030, new_AGEMA_signal_25027}), .clk (clk), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({new_AGEMA_signal_8018, new_AGEMA_signal_8017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7837, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_25042, new_AGEMA_signal_25039, new_AGEMA_signal_25036}), .clk (clk), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_25051, new_AGEMA_signal_25048, new_AGEMA_signal_25045}), .clk (clk), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_25060, new_AGEMA_signal_25057, new_AGEMA_signal_25054}), .clk (clk), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_25069, new_AGEMA_signal_25066, new_AGEMA_signal_25063}), .clk (clk), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_8006, new_AGEMA_signal_8005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_8486, new_AGEMA_signal_8485, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_8960, new_AGEMA_signal_8959, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_8480, new_AGEMA_signal_8479, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_8018, new_AGEMA_signal_8017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_8492, new_AGEMA_signal_8491, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_8972, new_AGEMA_signal_8971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_8966, new_AGEMA_signal_8965, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_9374, new_AGEMA_signal_9373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_8972, new_AGEMA_signal_8971, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_9362, new_AGEMA_signal_9361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_8498, new_AGEMA_signal_8497, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_9368, new_AGEMA_signal_9367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_10166, new_AGEMA_signal_10165, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_10172, new_AGEMA_signal_10171, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_10178, new_AGEMA_signal_10177, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_9374, new_AGEMA_signal_9373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_25078, new_AGEMA_signal_25075, new_AGEMA_signal_25072}), .clk (clk), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_25087, new_AGEMA_signal_25084, new_AGEMA_signal_25081}), .clk (clk), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({new_AGEMA_signal_8030, new_AGEMA_signal_8029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_23371, new_AGEMA_signal_23367, new_AGEMA_signal_23363}), .clk (clk), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_25096, new_AGEMA_signal_25093, new_AGEMA_signal_25090}), .clk (clk), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_25105, new_AGEMA_signal_25102, new_AGEMA_signal_25099}), .clk (clk), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_25114, new_AGEMA_signal_25111, new_AGEMA_signal_25108}), .clk (clk), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_25123, new_AGEMA_signal_25120, new_AGEMA_signal_25117}), .clk (clk), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_25132, new_AGEMA_signal_25129, new_AGEMA_signal_25126}), .clk (clk), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_25141, new_AGEMA_signal_25138, new_AGEMA_signal_25135}), .clk (clk), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({new_AGEMA_signal_8510, new_AGEMA_signal_8509, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_25150, new_AGEMA_signal_25147, new_AGEMA_signal_25144}), .clk (clk), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_25159, new_AGEMA_signal_25156, new_AGEMA_signal_25153}), .clk (clk), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7849, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_25168, new_AGEMA_signal_25165, new_AGEMA_signal_25162}), .clk (clk), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_25177, new_AGEMA_signal_25174, new_AGEMA_signal_25171}), .clk (clk), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_25186, new_AGEMA_signal_25183, new_AGEMA_signal_25180}), .clk (clk), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({new_AGEMA_signal_8042, new_AGEMA_signal_8041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_25195, new_AGEMA_signal_25192, new_AGEMA_signal_25189}), .clk (clk), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_8024, new_AGEMA_signal_8023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_25204, new_AGEMA_signal_25201, new_AGEMA_signal_25198}), .clk (clk), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_25213, new_AGEMA_signal_25210, new_AGEMA_signal_25207}), .clk (clk), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_25222, new_AGEMA_signal_25219, new_AGEMA_signal_25216}), .clk (clk), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_8030, new_AGEMA_signal_8029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_8510, new_AGEMA_signal_8509, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_8504, new_AGEMA_signal_8503, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_8042, new_AGEMA_signal_8041, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_8978, new_AGEMA_signal_8977, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_8036, new_AGEMA_signal_8035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_8516, new_AGEMA_signal_8515, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_8990, new_AGEMA_signal_8989, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_8996, new_AGEMA_signal_8995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_8984, new_AGEMA_signal_8983, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_8996, new_AGEMA_signal_8995, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_9392, new_AGEMA_signal_9391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_9380, new_AGEMA_signal_9379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_8522, new_AGEMA_signal_8521, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_8990, new_AGEMA_signal_8989, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_10184, new_AGEMA_signal_10183, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_10190, new_AGEMA_signal_10189, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_9392, new_AGEMA_signal_9391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_25231, new_AGEMA_signal_25228, new_AGEMA_signal_25225}), .clk (clk), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_25240, new_AGEMA_signal_25237, new_AGEMA_signal_25234}), .clk (clk), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({new_AGEMA_signal_8054, new_AGEMA_signal_8053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_24847, new_AGEMA_signal_24843, new_AGEMA_signal_24839}), .clk (clk), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_25249, new_AGEMA_signal_25246, new_AGEMA_signal_25243}), .clk (clk), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_25258, new_AGEMA_signal_25255, new_AGEMA_signal_25252}), .clk (clk), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_25267, new_AGEMA_signal_25264, new_AGEMA_signal_25261}), .clk (clk), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_25276, new_AGEMA_signal_25273, new_AGEMA_signal_25270}), .clk (clk), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_25285, new_AGEMA_signal_25282, new_AGEMA_signal_25279}), .clk (clk), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_25294, new_AGEMA_signal_25291, new_AGEMA_signal_25288}), .clk (clk), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({new_AGEMA_signal_8534, new_AGEMA_signal_8533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_25303, new_AGEMA_signal_25300, new_AGEMA_signal_25297}), .clk (clk), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_25312, new_AGEMA_signal_25309, new_AGEMA_signal_25306}), .clk (clk), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_25321, new_AGEMA_signal_25318, new_AGEMA_signal_25315}), .clk (clk), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_25330, new_AGEMA_signal_25327, new_AGEMA_signal_25324}), .clk (clk), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_7856, new_AGEMA_signal_7855, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_25339, new_AGEMA_signal_25336, new_AGEMA_signal_25333}), .clk (clk), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({new_AGEMA_signal_8066, new_AGEMA_signal_8065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_25348, new_AGEMA_signal_25345, new_AGEMA_signal_25342}), .clk (clk), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_25357, new_AGEMA_signal_25354, new_AGEMA_signal_25351}), .clk (clk), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_25366, new_AGEMA_signal_25363, new_AGEMA_signal_25360}), .clk (clk), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_25375, new_AGEMA_signal_25372, new_AGEMA_signal_25369}), .clk (clk), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_8054, new_AGEMA_signal_8053, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_8534, new_AGEMA_signal_8533, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9008, new_AGEMA_signal_9007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_9008, new_AGEMA_signal_9007, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_8528, new_AGEMA_signal_8527, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_8066, new_AGEMA_signal_8065, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_8060, new_AGEMA_signal_8059, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_8540, new_AGEMA_signal_8539, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9014, new_AGEMA_signal_9013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9001, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_9410, new_AGEMA_signal_9409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_9398, new_AGEMA_signal_9397, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_8546, new_AGEMA_signal_8545, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_9404, new_AGEMA_signal_9403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_9014, new_AGEMA_signal_9013, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_10196, new_AGEMA_signal_10195, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_10202, new_AGEMA_signal_10201, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_9410, new_AGEMA_signal_9409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_25384, new_AGEMA_signal_25381, new_AGEMA_signal_25378}), .clk (clk), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_25393, new_AGEMA_signal_25390, new_AGEMA_signal_25387}), .clk (clk), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({new_AGEMA_signal_8078, new_AGEMA_signal_8077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_23923, new_AGEMA_signal_23919, new_AGEMA_signal_23915}), .clk (clk), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_25402, new_AGEMA_signal_25399, new_AGEMA_signal_25396}), .clk (clk), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_25411, new_AGEMA_signal_25408, new_AGEMA_signal_25405}), .clk (clk), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_25420, new_AGEMA_signal_25417, new_AGEMA_signal_25414}), .clk (clk), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_25429, new_AGEMA_signal_25426, new_AGEMA_signal_25423}), .clk (clk), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_25438, new_AGEMA_signal_25435, new_AGEMA_signal_25432}), .clk (clk), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_25447, new_AGEMA_signal_25444, new_AGEMA_signal_25441}), .clk (clk), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({new_AGEMA_signal_8558, new_AGEMA_signal_8557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_25456, new_AGEMA_signal_25453, new_AGEMA_signal_25450}), .clk (clk), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_7868, new_AGEMA_signal_7867, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_25465, new_AGEMA_signal_25462, new_AGEMA_signal_25459}), .clk (clk), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_25474, new_AGEMA_signal_25471, new_AGEMA_signal_25468}), .clk (clk), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_25483, new_AGEMA_signal_25480, new_AGEMA_signal_25477}), .clk (clk), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_25492, new_AGEMA_signal_25489, new_AGEMA_signal_25486}), .clk (clk), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({new_AGEMA_signal_8090, new_AGEMA_signal_8089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7861, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_25501, new_AGEMA_signal_25498, new_AGEMA_signal_25495}), .clk (clk), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8071, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_25510, new_AGEMA_signal_25507, new_AGEMA_signal_25504}), .clk (clk), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_25519, new_AGEMA_signal_25516, new_AGEMA_signal_25513}), .clk (clk), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_25528, new_AGEMA_signal_25525, new_AGEMA_signal_25522}), .clk (clk), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_8078, new_AGEMA_signal_8077, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_8558, new_AGEMA_signal_8557, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_9020, new_AGEMA_signal_9019, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_8552, new_AGEMA_signal_8551, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_8090, new_AGEMA_signal_8089, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_8564, new_AGEMA_signal_8563, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9032, new_AGEMA_signal_9031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_9026, new_AGEMA_signal_9025, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_9428, new_AGEMA_signal_9427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_9032, new_AGEMA_signal_9031, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_9416, new_AGEMA_signal_9415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_8570, new_AGEMA_signal_8569, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_9422, new_AGEMA_signal_9421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_10208, new_AGEMA_signal_10207, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_10214, new_AGEMA_signal_10213, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_10220, new_AGEMA_signal_10219, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_9428, new_AGEMA_signal_9427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, KeyExpansionIns_tmp[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_17655), .Q (new_AGEMA_signal_17656) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_17659), .Q (new_AGEMA_signal_17660) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_17663), .Q (new_AGEMA_signal_17664) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_17667), .Q (new_AGEMA_signal_17668) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_17671), .Q (new_AGEMA_signal_17672) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_17675), .Q (new_AGEMA_signal_17676) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_17679), .Q (new_AGEMA_signal_17680) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_17683), .Q (new_AGEMA_signal_17684) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_17687), .Q (new_AGEMA_signal_17688) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_17691), .Q (new_AGEMA_signal_17692) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_17695), .Q (new_AGEMA_signal_17696) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_17699), .Q (new_AGEMA_signal_17700) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_17703), .Q (new_AGEMA_signal_17704) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_17707), .Q (new_AGEMA_signal_17708) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_17711), .Q (new_AGEMA_signal_17712) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_17715), .Q (new_AGEMA_signal_17716) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_17719), .Q (new_AGEMA_signal_17720) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_17723), .Q (new_AGEMA_signal_17724) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_17727), .Q (new_AGEMA_signal_17728) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_17731), .Q (new_AGEMA_signal_17732) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_17735), .Q (new_AGEMA_signal_17736) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_17739), .Q (new_AGEMA_signal_17740) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_17743), .Q (new_AGEMA_signal_17744) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_17747), .Q (new_AGEMA_signal_17748) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_17751), .Q (new_AGEMA_signal_17752) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_17755), .Q (new_AGEMA_signal_17756) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_17759), .Q (new_AGEMA_signal_17760) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_17763), .Q (new_AGEMA_signal_17764) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_17767), .Q (new_AGEMA_signal_17768) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_17771), .Q (new_AGEMA_signal_17772) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_17775), .Q (new_AGEMA_signal_17776) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_17779), .Q (new_AGEMA_signal_17780) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_17783), .Q (new_AGEMA_signal_17784) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_17787), .Q (new_AGEMA_signal_17788) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_17791), .Q (new_AGEMA_signal_17792) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_17795), .Q (new_AGEMA_signal_17796) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_17799), .Q (new_AGEMA_signal_17800) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_17803), .Q (new_AGEMA_signal_17804) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_17807), .Q (new_AGEMA_signal_17808) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_17811), .Q (new_AGEMA_signal_17812) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_17815), .Q (new_AGEMA_signal_17816) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_17819), .Q (new_AGEMA_signal_17820) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_17823), .Q (new_AGEMA_signal_17824) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_17827), .Q (new_AGEMA_signal_17828) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_17831), .Q (new_AGEMA_signal_17832) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_17835), .Q (new_AGEMA_signal_17836) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_17839), .Q (new_AGEMA_signal_17840) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_17843), .Q (new_AGEMA_signal_17844) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_17847), .Q (new_AGEMA_signal_17848) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_17851), .Q (new_AGEMA_signal_17852) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_17855), .Q (new_AGEMA_signal_17856) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_17859), .Q (new_AGEMA_signal_17860) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_17863), .Q (new_AGEMA_signal_17864) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_17867), .Q (new_AGEMA_signal_17868) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_17871), .Q (new_AGEMA_signal_17872) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_17875), .Q (new_AGEMA_signal_17876) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_17879), .Q (new_AGEMA_signal_17880) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_17883), .Q (new_AGEMA_signal_17884) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_17887), .Q (new_AGEMA_signal_17888) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_17891), .Q (new_AGEMA_signal_17892) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_17895), .Q (new_AGEMA_signal_17896) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_17899), .Q (new_AGEMA_signal_17900) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_17903), .Q (new_AGEMA_signal_17904) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_17907), .Q (new_AGEMA_signal_17908) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_17911), .Q (new_AGEMA_signal_17912) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_17915), .Q (new_AGEMA_signal_17916) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_17919), .Q (new_AGEMA_signal_17920) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_17923), .Q (new_AGEMA_signal_17924) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_17927), .Q (new_AGEMA_signal_17928) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_17931), .Q (new_AGEMA_signal_17932) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_17935), .Q (new_AGEMA_signal_17936) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_17939), .Q (new_AGEMA_signal_17940) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_17943), .Q (new_AGEMA_signal_17944) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_17947), .Q (new_AGEMA_signal_17948) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_17951), .Q (new_AGEMA_signal_17952) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_17955), .Q (new_AGEMA_signal_17956) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_17959), .Q (new_AGEMA_signal_17960) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_17963), .Q (new_AGEMA_signal_17964) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_17967), .Q (new_AGEMA_signal_17968) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_17971), .Q (new_AGEMA_signal_17972) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_17975), .Q (new_AGEMA_signal_17976) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_17979), .Q (new_AGEMA_signal_17980) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_17983), .Q (new_AGEMA_signal_17984) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_17987), .Q (new_AGEMA_signal_17988) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_17991), .Q (new_AGEMA_signal_17992) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_17995), .Q (new_AGEMA_signal_17996) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_17999), .Q (new_AGEMA_signal_18000) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_18003), .Q (new_AGEMA_signal_18004) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_18007), .Q (new_AGEMA_signal_18008) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_18011), .Q (new_AGEMA_signal_18012) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_18015), .Q (new_AGEMA_signal_18016) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_18019), .Q (new_AGEMA_signal_18020) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_18023), .Q (new_AGEMA_signal_18024) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_18027), .Q (new_AGEMA_signal_18028) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_18031), .Q (new_AGEMA_signal_18032) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_18035), .Q (new_AGEMA_signal_18036) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_18039), .Q (new_AGEMA_signal_18040) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_18043), .Q (new_AGEMA_signal_18044) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_18047), .Q (new_AGEMA_signal_18048) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_18051), .Q (new_AGEMA_signal_18052) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_18055), .Q (new_AGEMA_signal_18056) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_18059), .Q (new_AGEMA_signal_18060) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_18063), .Q (new_AGEMA_signal_18064) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_18067), .Q (new_AGEMA_signal_18068) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_18071), .Q (new_AGEMA_signal_18072) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_18075), .Q (new_AGEMA_signal_18076) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_18079), .Q (new_AGEMA_signal_18080) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_18083), .Q (new_AGEMA_signal_18084) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_18087), .Q (new_AGEMA_signal_18088) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_18091), .Q (new_AGEMA_signal_18092) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_18095), .Q (new_AGEMA_signal_18096) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_18099), .Q (new_AGEMA_signal_18100) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_18103), .Q (new_AGEMA_signal_18104) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_18107), .Q (new_AGEMA_signal_18108) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_18111), .Q (new_AGEMA_signal_18112) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_18115), .Q (new_AGEMA_signal_18116) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_18119), .Q (new_AGEMA_signal_18120) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_18123), .Q (new_AGEMA_signal_18124) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_18127), .Q (new_AGEMA_signal_18128) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_18131), .Q (new_AGEMA_signal_18132) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_18135), .Q (new_AGEMA_signal_18136) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_18139), .Q (new_AGEMA_signal_18140) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_18143), .Q (new_AGEMA_signal_18144) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_18147), .Q (new_AGEMA_signal_18148) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_18151), .Q (new_AGEMA_signal_18152) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_18155), .Q (new_AGEMA_signal_18156) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_18159), .Q (new_AGEMA_signal_18160) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_18163), .Q (new_AGEMA_signal_18164) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_18167), .Q (new_AGEMA_signal_18168) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_18171), .Q (new_AGEMA_signal_18172) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_18175), .Q (new_AGEMA_signal_18176) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_18179), .Q (new_AGEMA_signal_18180) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_18183), .Q (new_AGEMA_signal_18184) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_18187), .Q (new_AGEMA_signal_18188) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_18191), .Q (new_AGEMA_signal_18192) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_18195), .Q (new_AGEMA_signal_18196) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_18199), .Q (new_AGEMA_signal_18200) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_18203), .Q (new_AGEMA_signal_18204) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_18207), .Q (new_AGEMA_signal_18208) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_18211), .Q (new_AGEMA_signal_18212) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_18215), .Q (new_AGEMA_signal_18216) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_18219), .Q (new_AGEMA_signal_18220) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_18223), .Q (new_AGEMA_signal_18224) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_18227), .Q (new_AGEMA_signal_18228) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_18231), .Q (new_AGEMA_signal_18232) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_18235), .Q (new_AGEMA_signal_18236) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_18239), .Q (new_AGEMA_signal_18240) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_18243), .Q (new_AGEMA_signal_18244) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_18247), .Q (new_AGEMA_signal_18248) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_18251), .Q (new_AGEMA_signal_18252) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_18255), .Q (new_AGEMA_signal_18256) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_18259), .Q (new_AGEMA_signal_18260) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_18263), .Q (new_AGEMA_signal_18264) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_18267), .Q (new_AGEMA_signal_18268) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_18271), .Q (new_AGEMA_signal_18272) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_18275), .Q (new_AGEMA_signal_18276) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_18279), .Q (new_AGEMA_signal_18280) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_18283), .Q (new_AGEMA_signal_18284) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_18287), .Q (new_AGEMA_signal_18288) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_18291), .Q (new_AGEMA_signal_18292) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_18295), .Q (new_AGEMA_signal_18296) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_18299), .Q (new_AGEMA_signal_18300) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_18303), .Q (new_AGEMA_signal_18304) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_18307), .Q (new_AGEMA_signal_18308) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_18311), .Q (new_AGEMA_signal_18312) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_18315), .Q (new_AGEMA_signal_18316) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_18319), .Q (new_AGEMA_signal_18320) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_18323), .Q (new_AGEMA_signal_18324) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_18327), .Q (new_AGEMA_signal_18328) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_18331), .Q (new_AGEMA_signal_18332) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_18335), .Q (new_AGEMA_signal_18336) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_18339), .Q (new_AGEMA_signal_18340) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_18343), .Q (new_AGEMA_signal_18344) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_18347), .Q (new_AGEMA_signal_18348) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_18351), .Q (new_AGEMA_signal_18352) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_18355), .Q (new_AGEMA_signal_18356) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_18359), .Q (new_AGEMA_signal_18360) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_18363), .Q (new_AGEMA_signal_18364) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_18367), .Q (new_AGEMA_signal_18368) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_18371), .Q (new_AGEMA_signal_18372) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_18375), .Q (new_AGEMA_signal_18376) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_18379), .Q (new_AGEMA_signal_18380) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_18383), .Q (new_AGEMA_signal_18384) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_18387), .Q (new_AGEMA_signal_18388) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_18391), .Q (new_AGEMA_signal_18392) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_18395), .Q (new_AGEMA_signal_18396) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_18399), .Q (new_AGEMA_signal_18400) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_18403), .Q (new_AGEMA_signal_18404) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_18407), .Q (new_AGEMA_signal_18408) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_18411), .Q (new_AGEMA_signal_18412) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_18415), .Q (new_AGEMA_signal_18416) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_18419), .Q (new_AGEMA_signal_18420) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_18423), .Q (new_AGEMA_signal_18424) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_18427), .Q (new_AGEMA_signal_18428) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_18431), .Q (new_AGEMA_signal_18432) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_18435), .Q (new_AGEMA_signal_18436) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_18439), .Q (new_AGEMA_signal_18440) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_18443), .Q (new_AGEMA_signal_18444) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_18447), .Q (new_AGEMA_signal_18448) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_18451), .Q (new_AGEMA_signal_18452) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_18455), .Q (new_AGEMA_signal_18456) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_18459), .Q (new_AGEMA_signal_18460) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_18463), .Q (new_AGEMA_signal_18464) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_18467), .Q (new_AGEMA_signal_18468) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_18471), .Q (new_AGEMA_signal_18472) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_18475), .Q (new_AGEMA_signal_18476) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_18479), .Q (new_AGEMA_signal_18480) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_18483), .Q (new_AGEMA_signal_18484) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_18487), .Q (new_AGEMA_signal_18488) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_18491), .Q (new_AGEMA_signal_18492) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_18495), .Q (new_AGEMA_signal_18496) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_18499), .Q (new_AGEMA_signal_18500) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_18503), .Q (new_AGEMA_signal_18504) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_18507), .Q (new_AGEMA_signal_18508) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_18511), .Q (new_AGEMA_signal_18512) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_18515), .Q (new_AGEMA_signal_18516) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_18519), .Q (new_AGEMA_signal_18520) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_18523), .Q (new_AGEMA_signal_18524) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_18527), .Q (new_AGEMA_signal_18528) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_18531), .Q (new_AGEMA_signal_18532) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_18535), .Q (new_AGEMA_signal_18536) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_18539), .Q (new_AGEMA_signal_18540) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_18543), .Q (new_AGEMA_signal_18544) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_18547), .Q (new_AGEMA_signal_18548) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_18551), .Q (new_AGEMA_signal_18552) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_18555), .Q (new_AGEMA_signal_18556) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_18559), .Q (new_AGEMA_signal_18560) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_18563), .Q (new_AGEMA_signal_18564) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_18567), .Q (new_AGEMA_signal_18568) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_18571), .Q (new_AGEMA_signal_18572) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_18575), .Q (new_AGEMA_signal_18576) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_18579), .Q (new_AGEMA_signal_18580) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_18583), .Q (new_AGEMA_signal_18584) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_18587), .Q (new_AGEMA_signal_18588) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_18591), .Q (new_AGEMA_signal_18592) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_18595), .Q (new_AGEMA_signal_18596) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_18599), .Q (new_AGEMA_signal_18600) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_18603), .Q (new_AGEMA_signal_18604) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_18607), .Q (new_AGEMA_signal_18608) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_18611), .Q (new_AGEMA_signal_18612) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_18615), .Q (new_AGEMA_signal_18616) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_18619), .Q (new_AGEMA_signal_18620) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_18623), .Q (new_AGEMA_signal_18624) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_18627), .Q (new_AGEMA_signal_18628) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_18631), .Q (new_AGEMA_signal_18632) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_18635), .Q (new_AGEMA_signal_18636) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_18639), .Q (new_AGEMA_signal_18640) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_18643), .Q (new_AGEMA_signal_18644) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_18647), .Q (new_AGEMA_signal_18648) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_18651), .Q (new_AGEMA_signal_18652) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_18655), .Q (new_AGEMA_signal_18656) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_18659), .Q (new_AGEMA_signal_18660) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_18663), .Q (new_AGEMA_signal_18664) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_18667), .Q (new_AGEMA_signal_18668) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_18671), .Q (new_AGEMA_signal_18672) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_18675), .Q (new_AGEMA_signal_18676) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_18679), .Q (new_AGEMA_signal_18680) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_18683), .Q (new_AGEMA_signal_18684) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_18687), .Q (new_AGEMA_signal_18688) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_18691), .Q (new_AGEMA_signal_18692) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_18695), .Q (new_AGEMA_signal_18696) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_18699), .Q (new_AGEMA_signal_18700) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_18703), .Q (new_AGEMA_signal_18704) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_18707), .Q (new_AGEMA_signal_18708) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_18711), .Q (new_AGEMA_signal_18712) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_18715), .Q (new_AGEMA_signal_18716) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_18719), .Q (new_AGEMA_signal_18720) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_18723), .Q (new_AGEMA_signal_18724) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_18727), .Q (new_AGEMA_signal_18728) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_18731), .Q (new_AGEMA_signal_18732) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_18735), .Q (new_AGEMA_signal_18736) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_18739), .Q (new_AGEMA_signal_18740) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_18743), .Q (new_AGEMA_signal_18744) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_18747), .Q (new_AGEMA_signal_18748) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_18751), .Q (new_AGEMA_signal_18752) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_18755), .Q (new_AGEMA_signal_18756) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_18759), .Q (new_AGEMA_signal_18760) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_18763), .Q (new_AGEMA_signal_18764) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_18767), .Q (new_AGEMA_signal_18768) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_18771), .Q (new_AGEMA_signal_18772) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_18775), .Q (new_AGEMA_signal_18776) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_18779), .Q (new_AGEMA_signal_18780) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_18783), .Q (new_AGEMA_signal_18784) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_18787), .Q (new_AGEMA_signal_18788) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_18791), .Q (new_AGEMA_signal_18792) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_18795), .Q (new_AGEMA_signal_18796) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_18799), .Q (new_AGEMA_signal_18800) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_18803), .Q (new_AGEMA_signal_18804) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C (clk), .D (new_AGEMA_signal_18807), .Q (new_AGEMA_signal_18808) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_18811), .Q (new_AGEMA_signal_18812) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_18815), .Q (new_AGEMA_signal_18816) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_18819), .Q (new_AGEMA_signal_18820) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_18823), .Q (new_AGEMA_signal_18824) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_18827), .Q (new_AGEMA_signal_18828) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_18831), .Q (new_AGEMA_signal_18832) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_18835), .Q (new_AGEMA_signal_18836) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_18839), .Q (new_AGEMA_signal_18840) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_18843), .Q (new_AGEMA_signal_18844) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_18847), .Q (new_AGEMA_signal_18848) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_18851), .Q (new_AGEMA_signal_18852) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_18855), .Q (new_AGEMA_signal_18856) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_18859), .Q (new_AGEMA_signal_18860) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_18863), .Q (new_AGEMA_signal_18864) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_18867), .Q (new_AGEMA_signal_18868) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_18871), .Q (new_AGEMA_signal_18872) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_18875), .Q (new_AGEMA_signal_18876) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_18879), .Q (new_AGEMA_signal_18880) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_18883), .Q (new_AGEMA_signal_18884) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_18887), .Q (new_AGEMA_signal_18888) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_18891), .Q (new_AGEMA_signal_18892) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_18895), .Q (new_AGEMA_signal_18896) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_18899), .Q (new_AGEMA_signal_18900) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_18903), .Q (new_AGEMA_signal_18904) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_18907), .Q (new_AGEMA_signal_18908) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_18911), .Q (new_AGEMA_signal_18912) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C (clk), .D (new_AGEMA_signal_18915), .Q (new_AGEMA_signal_18916) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_18919), .Q (new_AGEMA_signal_18920) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_18923), .Q (new_AGEMA_signal_18924) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_18927), .Q (new_AGEMA_signal_18928) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_18931), .Q (new_AGEMA_signal_18932) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_18935), .Q (new_AGEMA_signal_18936) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_18939), .Q (new_AGEMA_signal_18940) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_18943), .Q (new_AGEMA_signal_18944) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_18947), .Q (new_AGEMA_signal_18948) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_18951), .Q (new_AGEMA_signal_18952) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_18955), .Q (new_AGEMA_signal_18956) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_18959), .Q (new_AGEMA_signal_18960) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_18963), .Q (new_AGEMA_signal_18964) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_18967), .Q (new_AGEMA_signal_18968) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_18971), .Q (new_AGEMA_signal_18972) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_18975), .Q (new_AGEMA_signal_18976) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_18979), .Q (new_AGEMA_signal_18980) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_18983), .Q (new_AGEMA_signal_18984) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_18987), .Q (new_AGEMA_signal_18988) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_18991), .Q (new_AGEMA_signal_18992) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_18995), .Q (new_AGEMA_signal_18996) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_18999), .Q (new_AGEMA_signal_19000) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_19003), .Q (new_AGEMA_signal_19004) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_19007), .Q (new_AGEMA_signal_19008) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_19011), .Q (new_AGEMA_signal_19012) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_19015), .Q (new_AGEMA_signal_19016) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_19019), .Q (new_AGEMA_signal_19020) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C (clk), .D (new_AGEMA_signal_19023), .Q (new_AGEMA_signal_19024) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_19027), .Q (new_AGEMA_signal_19028) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_19031), .Q (new_AGEMA_signal_19032) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_19035), .Q (new_AGEMA_signal_19036) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_19039), .Q (new_AGEMA_signal_19040) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_19043), .Q (new_AGEMA_signal_19044) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_19047), .Q (new_AGEMA_signal_19048) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_19051), .Q (new_AGEMA_signal_19052) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_19055), .Q (new_AGEMA_signal_19056) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_19059), .Q (new_AGEMA_signal_19060) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_19063), .Q (new_AGEMA_signal_19064) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_19067), .Q (new_AGEMA_signal_19068) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_19071), .Q (new_AGEMA_signal_19072) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_19075), .Q (new_AGEMA_signal_19076) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_19079), .Q (new_AGEMA_signal_19080) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_19083), .Q (new_AGEMA_signal_19084) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_19087), .Q (new_AGEMA_signal_19088) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_19091), .Q (new_AGEMA_signal_19092) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_19095), .Q (new_AGEMA_signal_19096) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_19099), .Q (new_AGEMA_signal_19100) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_19103), .Q (new_AGEMA_signal_19104) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_19107), .Q (new_AGEMA_signal_19108) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_19111), .Q (new_AGEMA_signal_19112) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_19115), .Q (new_AGEMA_signal_19116) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_19119), .Q (new_AGEMA_signal_19120) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_19123), .Q (new_AGEMA_signal_19124) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_19127), .Q (new_AGEMA_signal_19128) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C (clk), .D (new_AGEMA_signal_19131), .Q (new_AGEMA_signal_19132) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_19135), .Q (new_AGEMA_signal_19136) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_19139), .Q (new_AGEMA_signal_19140) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_19143), .Q (new_AGEMA_signal_19144) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_19147), .Q (new_AGEMA_signal_19148) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_19151), .Q (new_AGEMA_signal_19152) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_19155), .Q (new_AGEMA_signal_19156) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_19159), .Q (new_AGEMA_signal_19160) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_19163), .Q (new_AGEMA_signal_19164) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_19167), .Q (new_AGEMA_signal_19168) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_19171), .Q (new_AGEMA_signal_19172) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_19175), .Q (new_AGEMA_signal_19176) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_19179), .Q (new_AGEMA_signal_19180) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_19183), .Q (new_AGEMA_signal_19184) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_19187), .Q (new_AGEMA_signal_19188) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_19191), .Q (new_AGEMA_signal_19192) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_19195), .Q (new_AGEMA_signal_19196) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_19199), .Q (new_AGEMA_signal_19200) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_19203), .Q (new_AGEMA_signal_19204) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_19207), .Q (new_AGEMA_signal_19208) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_19211), .Q (new_AGEMA_signal_19212) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_19215), .Q (new_AGEMA_signal_19216) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_19219), .Q (new_AGEMA_signal_19220) ) ;
    buf_clk new_AGEMA_reg_buffer_9092 ( .C (clk), .D (new_AGEMA_signal_21815), .Q (new_AGEMA_signal_21816) ) ;
    buf_clk new_AGEMA_reg_buffer_9096 ( .C (clk), .D (new_AGEMA_signal_21819), .Q (new_AGEMA_signal_21820) ) ;
    buf_clk new_AGEMA_reg_buffer_9100 ( .C (clk), .D (new_AGEMA_signal_21823), .Q (new_AGEMA_signal_21824) ) ;
    buf_clk new_AGEMA_reg_buffer_9104 ( .C (clk), .D (new_AGEMA_signal_21827), .Q (new_AGEMA_signal_21828) ) ;
    buf_clk new_AGEMA_reg_buffer_9108 ( .C (clk), .D (new_AGEMA_signal_21831), .Q (new_AGEMA_signal_21832) ) ;
    buf_clk new_AGEMA_reg_buffer_9112 ( .C (clk), .D (new_AGEMA_signal_21835), .Q (new_AGEMA_signal_21836) ) ;
    buf_clk new_AGEMA_reg_buffer_9116 ( .C (clk), .D (new_AGEMA_signal_21839), .Q (new_AGEMA_signal_21840) ) ;
    buf_clk new_AGEMA_reg_buffer_9120 ( .C (clk), .D (new_AGEMA_signal_21843), .Q (new_AGEMA_signal_21844) ) ;
    buf_clk new_AGEMA_reg_buffer_9124 ( .C (clk), .D (new_AGEMA_signal_21847), .Q (new_AGEMA_signal_21848) ) ;
    buf_clk new_AGEMA_reg_buffer_9128 ( .C (clk), .D (new_AGEMA_signal_21851), .Q (new_AGEMA_signal_21852) ) ;
    buf_clk new_AGEMA_reg_buffer_9132 ( .C (clk), .D (new_AGEMA_signal_21855), .Q (new_AGEMA_signal_21856) ) ;
    buf_clk new_AGEMA_reg_buffer_9136 ( .C (clk), .D (new_AGEMA_signal_21859), .Q (new_AGEMA_signal_21860) ) ;
    buf_clk new_AGEMA_reg_buffer_9140 ( .C (clk), .D (new_AGEMA_signal_21863), .Q (new_AGEMA_signal_21864) ) ;
    buf_clk new_AGEMA_reg_buffer_9144 ( .C (clk), .D (new_AGEMA_signal_21867), .Q (new_AGEMA_signal_21868) ) ;
    buf_clk new_AGEMA_reg_buffer_9148 ( .C (clk), .D (new_AGEMA_signal_21871), .Q (new_AGEMA_signal_21872) ) ;
    buf_clk new_AGEMA_reg_buffer_9152 ( .C (clk), .D (new_AGEMA_signal_21875), .Q (new_AGEMA_signal_21876) ) ;
    buf_clk new_AGEMA_reg_buffer_9156 ( .C (clk), .D (new_AGEMA_signal_21879), .Q (new_AGEMA_signal_21880) ) ;
    buf_clk new_AGEMA_reg_buffer_9160 ( .C (clk), .D (new_AGEMA_signal_21883), .Q (new_AGEMA_signal_21884) ) ;
    buf_clk new_AGEMA_reg_buffer_9164 ( .C (clk), .D (new_AGEMA_signal_21887), .Q (new_AGEMA_signal_21888) ) ;
    buf_clk new_AGEMA_reg_buffer_9168 ( .C (clk), .D (new_AGEMA_signal_21891), .Q (new_AGEMA_signal_21892) ) ;
    buf_clk new_AGEMA_reg_buffer_9172 ( .C (clk), .D (new_AGEMA_signal_21895), .Q (new_AGEMA_signal_21896) ) ;
    buf_clk new_AGEMA_reg_buffer_9176 ( .C (clk), .D (new_AGEMA_signal_21899), .Q (new_AGEMA_signal_21900) ) ;
    buf_clk new_AGEMA_reg_buffer_9180 ( .C (clk), .D (new_AGEMA_signal_21903), .Q (new_AGEMA_signal_21904) ) ;
    buf_clk new_AGEMA_reg_buffer_9184 ( .C (clk), .D (new_AGEMA_signal_21907), .Q (new_AGEMA_signal_21908) ) ;
    buf_clk new_AGEMA_reg_buffer_9188 ( .C (clk), .D (new_AGEMA_signal_21911), .Q (new_AGEMA_signal_21912) ) ;
    buf_clk new_AGEMA_reg_buffer_9192 ( .C (clk), .D (new_AGEMA_signal_21915), .Q (new_AGEMA_signal_21916) ) ;
    buf_clk new_AGEMA_reg_buffer_9196 ( .C (clk), .D (new_AGEMA_signal_21919), .Q (new_AGEMA_signal_21920) ) ;
    buf_clk new_AGEMA_reg_buffer_9200 ( .C (clk), .D (new_AGEMA_signal_21923), .Q (new_AGEMA_signal_21924) ) ;
    buf_clk new_AGEMA_reg_buffer_9204 ( .C (clk), .D (new_AGEMA_signal_21927), .Q (new_AGEMA_signal_21928) ) ;
    buf_clk new_AGEMA_reg_buffer_9208 ( .C (clk), .D (new_AGEMA_signal_21931), .Q (new_AGEMA_signal_21932) ) ;
    buf_clk new_AGEMA_reg_buffer_9212 ( .C (clk), .D (new_AGEMA_signal_21935), .Q (new_AGEMA_signal_21936) ) ;
    buf_clk new_AGEMA_reg_buffer_9216 ( .C (clk), .D (new_AGEMA_signal_21939), .Q (new_AGEMA_signal_21940) ) ;
    buf_clk new_AGEMA_reg_buffer_9220 ( .C (clk), .D (new_AGEMA_signal_21943), .Q (new_AGEMA_signal_21944) ) ;
    buf_clk new_AGEMA_reg_buffer_9224 ( .C (clk), .D (new_AGEMA_signal_21947), .Q (new_AGEMA_signal_21948) ) ;
    buf_clk new_AGEMA_reg_buffer_9228 ( .C (clk), .D (new_AGEMA_signal_21951), .Q (new_AGEMA_signal_21952) ) ;
    buf_clk new_AGEMA_reg_buffer_9232 ( .C (clk), .D (new_AGEMA_signal_21955), .Q (new_AGEMA_signal_21956) ) ;
    buf_clk new_AGEMA_reg_buffer_9236 ( .C (clk), .D (new_AGEMA_signal_21959), .Q (new_AGEMA_signal_21960) ) ;
    buf_clk new_AGEMA_reg_buffer_9240 ( .C (clk), .D (new_AGEMA_signal_21963), .Q (new_AGEMA_signal_21964) ) ;
    buf_clk new_AGEMA_reg_buffer_9244 ( .C (clk), .D (new_AGEMA_signal_21967), .Q (new_AGEMA_signal_21968) ) ;
    buf_clk new_AGEMA_reg_buffer_9248 ( .C (clk), .D (new_AGEMA_signal_21971), .Q (new_AGEMA_signal_21972) ) ;
    buf_clk new_AGEMA_reg_buffer_9252 ( .C (clk), .D (new_AGEMA_signal_21975), .Q (new_AGEMA_signal_21976) ) ;
    buf_clk new_AGEMA_reg_buffer_9256 ( .C (clk), .D (new_AGEMA_signal_21979), .Q (new_AGEMA_signal_21980) ) ;
    buf_clk new_AGEMA_reg_buffer_9260 ( .C (clk), .D (new_AGEMA_signal_21983), .Q (new_AGEMA_signal_21984) ) ;
    buf_clk new_AGEMA_reg_buffer_9264 ( .C (clk), .D (new_AGEMA_signal_21987), .Q (new_AGEMA_signal_21988) ) ;
    buf_clk new_AGEMA_reg_buffer_9268 ( .C (clk), .D (new_AGEMA_signal_21991), .Q (new_AGEMA_signal_21992) ) ;
    buf_clk new_AGEMA_reg_buffer_9272 ( .C (clk), .D (new_AGEMA_signal_21995), .Q (new_AGEMA_signal_21996) ) ;
    buf_clk new_AGEMA_reg_buffer_9276 ( .C (clk), .D (new_AGEMA_signal_21999), .Q (new_AGEMA_signal_22000) ) ;
    buf_clk new_AGEMA_reg_buffer_9280 ( .C (clk), .D (new_AGEMA_signal_22003), .Q (new_AGEMA_signal_22004) ) ;
    buf_clk new_AGEMA_reg_buffer_9284 ( .C (clk), .D (new_AGEMA_signal_22007), .Q (new_AGEMA_signal_22008) ) ;
    buf_clk new_AGEMA_reg_buffer_9288 ( .C (clk), .D (new_AGEMA_signal_22011), .Q (new_AGEMA_signal_22012) ) ;
    buf_clk new_AGEMA_reg_buffer_9292 ( .C (clk), .D (new_AGEMA_signal_22015), .Q (new_AGEMA_signal_22016) ) ;
    buf_clk new_AGEMA_reg_buffer_9296 ( .C (clk), .D (new_AGEMA_signal_22019), .Q (new_AGEMA_signal_22020) ) ;
    buf_clk new_AGEMA_reg_buffer_9300 ( .C (clk), .D (new_AGEMA_signal_22023), .Q (new_AGEMA_signal_22024) ) ;
    buf_clk new_AGEMA_reg_buffer_9304 ( .C (clk), .D (new_AGEMA_signal_22027), .Q (new_AGEMA_signal_22028) ) ;
    buf_clk new_AGEMA_reg_buffer_9308 ( .C (clk), .D (new_AGEMA_signal_22031), .Q (new_AGEMA_signal_22032) ) ;
    buf_clk new_AGEMA_reg_buffer_9312 ( .C (clk), .D (new_AGEMA_signal_22035), .Q (new_AGEMA_signal_22036) ) ;
    buf_clk new_AGEMA_reg_buffer_9316 ( .C (clk), .D (new_AGEMA_signal_22039), .Q (new_AGEMA_signal_22040) ) ;
    buf_clk new_AGEMA_reg_buffer_9320 ( .C (clk), .D (new_AGEMA_signal_22043), .Q (new_AGEMA_signal_22044) ) ;
    buf_clk new_AGEMA_reg_buffer_9324 ( .C (clk), .D (new_AGEMA_signal_22047), .Q (new_AGEMA_signal_22048) ) ;
    buf_clk new_AGEMA_reg_buffer_9328 ( .C (clk), .D (new_AGEMA_signal_22051), .Q (new_AGEMA_signal_22052) ) ;
    buf_clk new_AGEMA_reg_buffer_9332 ( .C (clk), .D (new_AGEMA_signal_22055), .Q (new_AGEMA_signal_22056) ) ;
    buf_clk new_AGEMA_reg_buffer_9336 ( .C (clk), .D (new_AGEMA_signal_22059), .Q (new_AGEMA_signal_22060) ) ;
    buf_clk new_AGEMA_reg_buffer_9340 ( .C (clk), .D (new_AGEMA_signal_22063), .Q (new_AGEMA_signal_22064) ) ;
    buf_clk new_AGEMA_reg_buffer_9344 ( .C (clk), .D (new_AGEMA_signal_22067), .Q (new_AGEMA_signal_22068) ) ;
    buf_clk new_AGEMA_reg_buffer_9348 ( .C (clk), .D (new_AGEMA_signal_22071), .Q (new_AGEMA_signal_22072) ) ;
    buf_clk new_AGEMA_reg_buffer_9352 ( .C (clk), .D (new_AGEMA_signal_22075), .Q (new_AGEMA_signal_22076) ) ;
    buf_clk new_AGEMA_reg_buffer_9356 ( .C (clk), .D (new_AGEMA_signal_22079), .Q (new_AGEMA_signal_22080) ) ;
    buf_clk new_AGEMA_reg_buffer_9360 ( .C (clk), .D (new_AGEMA_signal_22083), .Q (new_AGEMA_signal_22084) ) ;
    buf_clk new_AGEMA_reg_buffer_9364 ( .C (clk), .D (new_AGEMA_signal_22087), .Q (new_AGEMA_signal_22088) ) ;
    buf_clk new_AGEMA_reg_buffer_9368 ( .C (clk), .D (new_AGEMA_signal_22091), .Q (new_AGEMA_signal_22092) ) ;
    buf_clk new_AGEMA_reg_buffer_9372 ( .C (clk), .D (new_AGEMA_signal_22095), .Q (new_AGEMA_signal_22096) ) ;
    buf_clk new_AGEMA_reg_buffer_9376 ( .C (clk), .D (new_AGEMA_signal_22099), .Q (new_AGEMA_signal_22100) ) ;
    buf_clk new_AGEMA_reg_buffer_9380 ( .C (clk), .D (new_AGEMA_signal_22103), .Q (new_AGEMA_signal_22104) ) ;
    buf_clk new_AGEMA_reg_buffer_9384 ( .C (clk), .D (new_AGEMA_signal_22107), .Q (new_AGEMA_signal_22108) ) ;
    buf_clk new_AGEMA_reg_buffer_9388 ( .C (clk), .D (new_AGEMA_signal_22111), .Q (new_AGEMA_signal_22112) ) ;
    buf_clk new_AGEMA_reg_buffer_9392 ( .C (clk), .D (new_AGEMA_signal_22115), .Q (new_AGEMA_signal_22116) ) ;
    buf_clk new_AGEMA_reg_buffer_9396 ( .C (clk), .D (new_AGEMA_signal_22119), .Q (new_AGEMA_signal_22120) ) ;
    buf_clk new_AGEMA_reg_buffer_9400 ( .C (clk), .D (new_AGEMA_signal_22123), .Q (new_AGEMA_signal_22124) ) ;
    buf_clk new_AGEMA_reg_buffer_9404 ( .C (clk), .D (new_AGEMA_signal_22127), .Q (new_AGEMA_signal_22128) ) ;
    buf_clk new_AGEMA_reg_buffer_9408 ( .C (clk), .D (new_AGEMA_signal_22131), .Q (new_AGEMA_signal_22132) ) ;
    buf_clk new_AGEMA_reg_buffer_9412 ( .C (clk), .D (new_AGEMA_signal_22135), .Q (new_AGEMA_signal_22136) ) ;
    buf_clk new_AGEMA_reg_buffer_9416 ( .C (clk), .D (new_AGEMA_signal_22139), .Q (new_AGEMA_signal_22140) ) ;
    buf_clk new_AGEMA_reg_buffer_9420 ( .C (clk), .D (new_AGEMA_signal_22143), .Q (new_AGEMA_signal_22144) ) ;
    buf_clk new_AGEMA_reg_buffer_9424 ( .C (clk), .D (new_AGEMA_signal_22147), .Q (new_AGEMA_signal_22148) ) ;
    buf_clk new_AGEMA_reg_buffer_9428 ( .C (clk), .D (new_AGEMA_signal_22151), .Q (new_AGEMA_signal_22152) ) ;
    buf_clk new_AGEMA_reg_buffer_9432 ( .C (clk), .D (new_AGEMA_signal_22155), .Q (new_AGEMA_signal_22156) ) ;
    buf_clk new_AGEMA_reg_buffer_9436 ( .C (clk), .D (new_AGEMA_signal_22159), .Q (new_AGEMA_signal_22160) ) ;
    buf_clk new_AGEMA_reg_buffer_9440 ( .C (clk), .D (new_AGEMA_signal_22163), .Q (new_AGEMA_signal_22164) ) ;
    buf_clk new_AGEMA_reg_buffer_9444 ( .C (clk), .D (new_AGEMA_signal_22167), .Q (new_AGEMA_signal_22168) ) ;
    buf_clk new_AGEMA_reg_buffer_9448 ( .C (clk), .D (new_AGEMA_signal_22171), .Q (new_AGEMA_signal_22172) ) ;
    buf_clk new_AGEMA_reg_buffer_9452 ( .C (clk), .D (new_AGEMA_signal_22175), .Q (new_AGEMA_signal_22176) ) ;
    buf_clk new_AGEMA_reg_buffer_9456 ( .C (clk), .D (new_AGEMA_signal_22179), .Q (new_AGEMA_signal_22180) ) ;
    buf_clk new_AGEMA_reg_buffer_9460 ( .C (clk), .D (new_AGEMA_signal_22183), .Q (new_AGEMA_signal_22184) ) ;
    buf_clk new_AGEMA_reg_buffer_9464 ( .C (clk), .D (new_AGEMA_signal_22187), .Q (new_AGEMA_signal_22188) ) ;
    buf_clk new_AGEMA_reg_buffer_9468 ( .C (clk), .D (new_AGEMA_signal_22191), .Q (new_AGEMA_signal_22192) ) ;
    buf_clk new_AGEMA_reg_buffer_9472 ( .C (clk), .D (new_AGEMA_signal_22195), .Q (new_AGEMA_signal_22196) ) ;
    buf_clk new_AGEMA_reg_buffer_9476 ( .C (clk), .D (new_AGEMA_signal_22199), .Q (new_AGEMA_signal_22200) ) ;
    buf_clk new_AGEMA_reg_buffer_9480 ( .C (clk), .D (new_AGEMA_signal_22203), .Q (new_AGEMA_signal_22204) ) ;
    buf_clk new_AGEMA_reg_buffer_9484 ( .C (clk), .D (new_AGEMA_signal_22207), .Q (new_AGEMA_signal_22208) ) ;
    buf_clk new_AGEMA_reg_buffer_9488 ( .C (clk), .D (new_AGEMA_signal_22211), .Q (new_AGEMA_signal_22212) ) ;
    buf_clk new_AGEMA_reg_buffer_9492 ( .C (clk), .D (new_AGEMA_signal_22215), .Q (new_AGEMA_signal_22216) ) ;
    buf_clk new_AGEMA_reg_buffer_9496 ( .C (clk), .D (new_AGEMA_signal_22219), .Q (new_AGEMA_signal_22220) ) ;
    buf_clk new_AGEMA_reg_buffer_9500 ( .C (clk), .D (new_AGEMA_signal_22223), .Q (new_AGEMA_signal_22224) ) ;
    buf_clk new_AGEMA_reg_buffer_9504 ( .C (clk), .D (new_AGEMA_signal_22227), .Q (new_AGEMA_signal_22228) ) ;
    buf_clk new_AGEMA_reg_buffer_9508 ( .C (clk), .D (new_AGEMA_signal_22231), .Q (new_AGEMA_signal_22232) ) ;
    buf_clk new_AGEMA_reg_buffer_9512 ( .C (clk), .D (new_AGEMA_signal_22235), .Q (new_AGEMA_signal_22236) ) ;
    buf_clk new_AGEMA_reg_buffer_9516 ( .C (clk), .D (new_AGEMA_signal_22239), .Q (new_AGEMA_signal_22240) ) ;
    buf_clk new_AGEMA_reg_buffer_9520 ( .C (clk), .D (new_AGEMA_signal_22243), .Q (new_AGEMA_signal_22244) ) ;
    buf_clk new_AGEMA_reg_buffer_9524 ( .C (clk), .D (new_AGEMA_signal_22247), .Q (new_AGEMA_signal_22248) ) ;
    buf_clk new_AGEMA_reg_buffer_9528 ( .C (clk), .D (new_AGEMA_signal_22251), .Q (new_AGEMA_signal_22252) ) ;
    buf_clk new_AGEMA_reg_buffer_9532 ( .C (clk), .D (new_AGEMA_signal_22255), .Q (new_AGEMA_signal_22256) ) ;
    buf_clk new_AGEMA_reg_buffer_9536 ( .C (clk), .D (new_AGEMA_signal_22259), .Q (new_AGEMA_signal_22260) ) ;
    buf_clk new_AGEMA_reg_buffer_9540 ( .C (clk), .D (new_AGEMA_signal_22263), .Q (new_AGEMA_signal_22264) ) ;
    buf_clk new_AGEMA_reg_buffer_9544 ( .C (clk), .D (new_AGEMA_signal_22267), .Q (new_AGEMA_signal_22268) ) ;
    buf_clk new_AGEMA_reg_buffer_9548 ( .C (clk), .D (new_AGEMA_signal_22271), .Q (new_AGEMA_signal_22272) ) ;
    buf_clk new_AGEMA_reg_buffer_9552 ( .C (clk), .D (new_AGEMA_signal_22275), .Q (new_AGEMA_signal_22276) ) ;
    buf_clk new_AGEMA_reg_buffer_9556 ( .C (clk), .D (new_AGEMA_signal_22279), .Q (new_AGEMA_signal_22280) ) ;
    buf_clk new_AGEMA_reg_buffer_9560 ( .C (clk), .D (new_AGEMA_signal_22283), .Q (new_AGEMA_signal_22284) ) ;
    buf_clk new_AGEMA_reg_buffer_9564 ( .C (clk), .D (new_AGEMA_signal_22287), .Q (new_AGEMA_signal_22288) ) ;
    buf_clk new_AGEMA_reg_buffer_9568 ( .C (clk), .D (new_AGEMA_signal_22291), .Q (new_AGEMA_signal_22292) ) ;
    buf_clk new_AGEMA_reg_buffer_9572 ( .C (clk), .D (new_AGEMA_signal_22295), .Q (new_AGEMA_signal_22296) ) ;
    buf_clk new_AGEMA_reg_buffer_9576 ( .C (clk), .D (new_AGEMA_signal_22299), .Q (new_AGEMA_signal_22300) ) ;
    buf_clk new_AGEMA_reg_buffer_9580 ( .C (clk), .D (new_AGEMA_signal_22303), .Q (new_AGEMA_signal_22304) ) ;
    buf_clk new_AGEMA_reg_buffer_9584 ( .C (clk), .D (new_AGEMA_signal_22307), .Q (new_AGEMA_signal_22308) ) ;
    buf_clk new_AGEMA_reg_buffer_9588 ( .C (clk), .D (new_AGEMA_signal_22311), .Q (new_AGEMA_signal_22312) ) ;
    buf_clk new_AGEMA_reg_buffer_9592 ( .C (clk), .D (new_AGEMA_signal_22315), .Q (new_AGEMA_signal_22316) ) ;
    buf_clk new_AGEMA_reg_buffer_9596 ( .C (clk), .D (new_AGEMA_signal_22319), .Q (new_AGEMA_signal_22320) ) ;
    buf_clk new_AGEMA_reg_buffer_9600 ( .C (clk), .D (new_AGEMA_signal_22323), .Q (new_AGEMA_signal_22324) ) ;
    buf_clk new_AGEMA_reg_buffer_9604 ( .C (clk), .D (new_AGEMA_signal_22327), .Q (new_AGEMA_signal_22328) ) ;
    buf_clk new_AGEMA_reg_buffer_9608 ( .C (clk), .D (new_AGEMA_signal_22331), .Q (new_AGEMA_signal_22332) ) ;
    buf_clk new_AGEMA_reg_buffer_9612 ( .C (clk), .D (new_AGEMA_signal_22335), .Q (new_AGEMA_signal_22336) ) ;
    buf_clk new_AGEMA_reg_buffer_9616 ( .C (clk), .D (new_AGEMA_signal_22339), .Q (new_AGEMA_signal_22340) ) ;
    buf_clk new_AGEMA_reg_buffer_9620 ( .C (clk), .D (new_AGEMA_signal_22343), .Q (new_AGEMA_signal_22344) ) ;
    buf_clk new_AGEMA_reg_buffer_9624 ( .C (clk), .D (new_AGEMA_signal_22347), .Q (new_AGEMA_signal_22348) ) ;
    buf_clk new_AGEMA_reg_buffer_9628 ( .C (clk), .D (new_AGEMA_signal_22351), .Q (new_AGEMA_signal_22352) ) ;
    buf_clk new_AGEMA_reg_buffer_9632 ( .C (clk), .D (new_AGEMA_signal_22355), .Q (new_AGEMA_signal_22356) ) ;
    buf_clk new_AGEMA_reg_buffer_9636 ( .C (clk), .D (new_AGEMA_signal_22359), .Q (new_AGEMA_signal_22360) ) ;
    buf_clk new_AGEMA_reg_buffer_9640 ( .C (clk), .D (new_AGEMA_signal_22363), .Q (new_AGEMA_signal_22364) ) ;
    buf_clk new_AGEMA_reg_buffer_9644 ( .C (clk), .D (new_AGEMA_signal_22367), .Q (new_AGEMA_signal_22368) ) ;
    buf_clk new_AGEMA_reg_buffer_9648 ( .C (clk), .D (new_AGEMA_signal_22371), .Q (new_AGEMA_signal_22372) ) ;
    buf_clk new_AGEMA_reg_buffer_9652 ( .C (clk), .D (new_AGEMA_signal_22375), .Q (new_AGEMA_signal_22376) ) ;
    buf_clk new_AGEMA_reg_buffer_9656 ( .C (clk), .D (new_AGEMA_signal_22379), .Q (new_AGEMA_signal_22380) ) ;
    buf_clk new_AGEMA_reg_buffer_9660 ( .C (clk), .D (new_AGEMA_signal_22383), .Q (new_AGEMA_signal_22384) ) ;
    buf_clk new_AGEMA_reg_buffer_9664 ( .C (clk), .D (new_AGEMA_signal_22387), .Q (new_AGEMA_signal_22388) ) ;
    buf_clk new_AGEMA_reg_buffer_9668 ( .C (clk), .D (new_AGEMA_signal_22391), .Q (new_AGEMA_signal_22392) ) ;
    buf_clk new_AGEMA_reg_buffer_9672 ( .C (clk), .D (new_AGEMA_signal_22395), .Q (new_AGEMA_signal_22396) ) ;
    buf_clk new_AGEMA_reg_buffer_9676 ( .C (clk), .D (new_AGEMA_signal_22399), .Q (new_AGEMA_signal_22400) ) ;
    buf_clk new_AGEMA_reg_buffer_9680 ( .C (clk), .D (new_AGEMA_signal_22403), .Q (new_AGEMA_signal_22404) ) ;
    buf_clk new_AGEMA_reg_buffer_9684 ( .C (clk), .D (new_AGEMA_signal_22407), .Q (new_AGEMA_signal_22408) ) ;
    buf_clk new_AGEMA_reg_buffer_9688 ( .C (clk), .D (new_AGEMA_signal_22411), .Q (new_AGEMA_signal_22412) ) ;
    buf_clk new_AGEMA_reg_buffer_9692 ( .C (clk), .D (new_AGEMA_signal_22415), .Q (new_AGEMA_signal_22416) ) ;
    buf_clk new_AGEMA_reg_buffer_9696 ( .C (clk), .D (new_AGEMA_signal_22419), .Q (new_AGEMA_signal_22420) ) ;
    buf_clk new_AGEMA_reg_buffer_9700 ( .C (clk), .D (new_AGEMA_signal_22423), .Q (new_AGEMA_signal_22424) ) ;
    buf_clk new_AGEMA_reg_buffer_9704 ( .C (clk), .D (new_AGEMA_signal_22427), .Q (new_AGEMA_signal_22428) ) ;
    buf_clk new_AGEMA_reg_buffer_9708 ( .C (clk), .D (new_AGEMA_signal_22431), .Q (new_AGEMA_signal_22432) ) ;
    buf_clk new_AGEMA_reg_buffer_9712 ( .C (clk), .D (new_AGEMA_signal_22435), .Q (new_AGEMA_signal_22436) ) ;
    buf_clk new_AGEMA_reg_buffer_9716 ( .C (clk), .D (new_AGEMA_signal_22439), .Q (new_AGEMA_signal_22440) ) ;
    buf_clk new_AGEMA_reg_buffer_9720 ( .C (clk), .D (new_AGEMA_signal_22443), .Q (new_AGEMA_signal_22444) ) ;
    buf_clk new_AGEMA_reg_buffer_9724 ( .C (clk), .D (new_AGEMA_signal_22447), .Q (new_AGEMA_signal_22448) ) ;
    buf_clk new_AGEMA_reg_buffer_9728 ( .C (clk), .D (new_AGEMA_signal_22451), .Q (new_AGEMA_signal_22452) ) ;
    buf_clk new_AGEMA_reg_buffer_9732 ( .C (clk), .D (new_AGEMA_signal_22455), .Q (new_AGEMA_signal_22456) ) ;
    buf_clk new_AGEMA_reg_buffer_9736 ( .C (clk), .D (new_AGEMA_signal_22459), .Q (new_AGEMA_signal_22460) ) ;
    buf_clk new_AGEMA_reg_buffer_9740 ( .C (clk), .D (new_AGEMA_signal_22463), .Q (new_AGEMA_signal_22464) ) ;
    buf_clk new_AGEMA_reg_buffer_9744 ( .C (clk), .D (new_AGEMA_signal_22467), .Q (new_AGEMA_signal_22468) ) ;
    buf_clk new_AGEMA_reg_buffer_9748 ( .C (clk), .D (new_AGEMA_signal_22471), .Q (new_AGEMA_signal_22472) ) ;
    buf_clk new_AGEMA_reg_buffer_9752 ( .C (clk), .D (new_AGEMA_signal_22475), .Q (new_AGEMA_signal_22476) ) ;
    buf_clk new_AGEMA_reg_buffer_9756 ( .C (clk), .D (new_AGEMA_signal_22479), .Q (new_AGEMA_signal_22480) ) ;
    buf_clk new_AGEMA_reg_buffer_9760 ( .C (clk), .D (new_AGEMA_signal_22483), .Q (new_AGEMA_signal_22484) ) ;
    buf_clk new_AGEMA_reg_buffer_9764 ( .C (clk), .D (new_AGEMA_signal_22487), .Q (new_AGEMA_signal_22488) ) ;
    buf_clk new_AGEMA_reg_buffer_9768 ( .C (clk), .D (new_AGEMA_signal_22491), .Q (new_AGEMA_signal_22492) ) ;
    buf_clk new_AGEMA_reg_buffer_9772 ( .C (clk), .D (new_AGEMA_signal_22495), .Q (new_AGEMA_signal_22496) ) ;
    buf_clk new_AGEMA_reg_buffer_9776 ( .C (clk), .D (new_AGEMA_signal_22499), .Q (new_AGEMA_signal_22500) ) ;
    buf_clk new_AGEMA_reg_buffer_9780 ( .C (clk), .D (new_AGEMA_signal_22503), .Q (new_AGEMA_signal_22504) ) ;
    buf_clk new_AGEMA_reg_buffer_9784 ( .C (clk), .D (new_AGEMA_signal_22507), .Q (new_AGEMA_signal_22508) ) ;
    buf_clk new_AGEMA_reg_buffer_9788 ( .C (clk), .D (new_AGEMA_signal_22511), .Q (new_AGEMA_signal_22512) ) ;
    buf_clk new_AGEMA_reg_buffer_9792 ( .C (clk), .D (new_AGEMA_signal_22515), .Q (new_AGEMA_signal_22516) ) ;
    buf_clk new_AGEMA_reg_buffer_9796 ( .C (clk), .D (new_AGEMA_signal_22519), .Q (new_AGEMA_signal_22520) ) ;
    buf_clk new_AGEMA_reg_buffer_9800 ( .C (clk), .D (new_AGEMA_signal_22523), .Q (new_AGEMA_signal_22524) ) ;
    buf_clk new_AGEMA_reg_buffer_9804 ( .C (clk), .D (new_AGEMA_signal_22527), .Q (new_AGEMA_signal_22528) ) ;
    buf_clk new_AGEMA_reg_buffer_9808 ( .C (clk), .D (new_AGEMA_signal_22531), .Q (new_AGEMA_signal_22532) ) ;
    buf_clk new_AGEMA_reg_buffer_9812 ( .C (clk), .D (new_AGEMA_signal_22535), .Q (new_AGEMA_signal_22536) ) ;
    buf_clk new_AGEMA_reg_buffer_9816 ( .C (clk), .D (new_AGEMA_signal_22539), .Q (new_AGEMA_signal_22540) ) ;
    buf_clk new_AGEMA_reg_buffer_9820 ( .C (clk), .D (new_AGEMA_signal_22543), .Q (new_AGEMA_signal_22544) ) ;
    buf_clk new_AGEMA_reg_buffer_9824 ( .C (clk), .D (new_AGEMA_signal_22547), .Q (new_AGEMA_signal_22548) ) ;
    buf_clk new_AGEMA_reg_buffer_9828 ( .C (clk), .D (new_AGEMA_signal_22551), .Q (new_AGEMA_signal_22552) ) ;
    buf_clk new_AGEMA_reg_buffer_9832 ( .C (clk), .D (new_AGEMA_signal_22555), .Q (new_AGEMA_signal_22556) ) ;
    buf_clk new_AGEMA_reg_buffer_9836 ( .C (clk), .D (new_AGEMA_signal_22559), .Q (new_AGEMA_signal_22560) ) ;
    buf_clk new_AGEMA_reg_buffer_9840 ( .C (clk), .D (new_AGEMA_signal_22563), .Q (new_AGEMA_signal_22564) ) ;
    buf_clk new_AGEMA_reg_buffer_9844 ( .C (clk), .D (new_AGEMA_signal_22567), .Q (new_AGEMA_signal_22568) ) ;
    buf_clk new_AGEMA_reg_buffer_9848 ( .C (clk), .D (new_AGEMA_signal_22571), .Q (new_AGEMA_signal_22572) ) ;
    buf_clk new_AGEMA_reg_buffer_9852 ( .C (clk), .D (new_AGEMA_signal_22575), .Q (new_AGEMA_signal_22576) ) ;
    buf_clk new_AGEMA_reg_buffer_9856 ( .C (clk), .D (new_AGEMA_signal_22579), .Q (new_AGEMA_signal_22580) ) ;
    buf_clk new_AGEMA_reg_buffer_9860 ( .C (clk), .D (new_AGEMA_signal_22583), .Q (new_AGEMA_signal_22584) ) ;
    buf_clk new_AGEMA_reg_buffer_9864 ( .C (clk), .D (new_AGEMA_signal_22587), .Q (new_AGEMA_signal_22588) ) ;
    buf_clk new_AGEMA_reg_buffer_9868 ( .C (clk), .D (new_AGEMA_signal_22591), .Q (new_AGEMA_signal_22592) ) ;
    buf_clk new_AGEMA_reg_buffer_9872 ( .C (clk), .D (new_AGEMA_signal_22595), .Q (new_AGEMA_signal_22596) ) ;
    buf_clk new_AGEMA_reg_buffer_9876 ( .C (clk), .D (new_AGEMA_signal_22599), .Q (new_AGEMA_signal_22600) ) ;
    buf_clk new_AGEMA_reg_buffer_9880 ( .C (clk), .D (new_AGEMA_signal_22603), .Q (new_AGEMA_signal_22604) ) ;
    buf_clk new_AGEMA_reg_buffer_9884 ( .C (clk), .D (new_AGEMA_signal_22607), .Q (new_AGEMA_signal_22608) ) ;
    buf_clk new_AGEMA_reg_buffer_9888 ( .C (clk), .D (new_AGEMA_signal_22611), .Q (new_AGEMA_signal_22612) ) ;
    buf_clk new_AGEMA_reg_buffer_9892 ( .C (clk), .D (new_AGEMA_signal_22615), .Q (new_AGEMA_signal_22616) ) ;
    buf_clk new_AGEMA_reg_buffer_9896 ( .C (clk), .D (new_AGEMA_signal_22619), .Q (new_AGEMA_signal_22620) ) ;
    buf_clk new_AGEMA_reg_buffer_9900 ( .C (clk), .D (new_AGEMA_signal_22623), .Q (new_AGEMA_signal_22624) ) ;
    buf_clk new_AGEMA_reg_buffer_9904 ( .C (clk), .D (new_AGEMA_signal_22627), .Q (new_AGEMA_signal_22628) ) ;
    buf_clk new_AGEMA_reg_buffer_9908 ( .C (clk), .D (new_AGEMA_signal_22631), .Q (new_AGEMA_signal_22632) ) ;
    buf_clk new_AGEMA_reg_buffer_9912 ( .C (clk), .D (new_AGEMA_signal_22635), .Q (new_AGEMA_signal_22636) ) ;
    buf_clk new_AGEMA_reg_buffer_9916 ( .C (clk), .D (new_AGEMA_signal_22639), .Q (new_AGEMA_signal_22640) ) ;
    buf_clk new_AGEMA_reg_buffer_9920 ( .C (clk), .D (new_AGEMA_signal_22643), .Q (new_AGEMA_signal_22644) ) ;
    buf_clk new_AGEMA_reg_buffer_9924 ( .C (clk), .D (new_AGEMA_signal_22647), .Q (new_AGEMA_signal_22648) ) ;
    buf_clk new_AGEMA_reg_buffer_9928 ( .C (clk), .D (new_AGEMA_signal_22651), .Q (new_AGEMA_signal_22652) ) ;
    buf_clk new_AGEMA_reg_buffer_9932 ( .C (clk), .D (new_AGEMA_signal_22655), .Q (new_AGEMA_signal_22656) ) ;
    buf_clk new_AGEMA_reg_buffer_9936 ( .C (clk), .D (new_AGEMA_signal_22659), .Q (new_AGEMA_signal_22660) ) ;
    buf_clk new_AGEMA_reg_buffer_9940 ( .C (clk), .D (new_AGEMA_signal_22663), .Q (new_AGEMA_signal_22664) ) ;
    buf_clk new_AGEMA_reg_buffer_9944 ( .C (clk), .D (new_AGEMA_signal_22667), .Q (new_AGEMA_signal_22668) ) ;
    buf_clk new_AGEMA_reg_buffer_9948 ( .C (clk), .D (new_AGEMA_signal_22671), .Q (new_AGEMA_signal_22672) ) ;
    buf_clk new_AGEMA_reg_buffer_9952 ( .C (clk), .D (new_AGEMA_signal_22675), .Q (new_AGEMA_signal_22676) ) ;
    buf_clk new_AGEMA_reg_buffer_9956 ( .C (clk), .D (new_AGEMA_signal_22679), .Q (new_AGEMA_signal_22680) ) ;
    buf_clk new_AGEMA_reg_buffer_9960 ( .C (clk), .D (new_AGEMA_signal_22683), .Q (new_AGEMA_signal_22684) ) ;
    buf_clk new_AGEMA_reg_buffer_9964 ( .C (clk), .D (new_AGEMA_signal_22687), .Q (new_AGEMA_signal_22688) ) ;
    buf_clk new_AGEMA_reg_buffer_9968 ( .C (clk), .D (new_AGEMA_signal_22691), .Q (new_AGEMA_signal_22692) ) ;
    buf_clk new_AGEMA_reg_buffer_9972 ( .C (clk), .D (new_AGEMA_signal_22695), .Q (new_AGEMA_signal_22696) ) ;
    buf_clk new_AGEMA_reg_buffer_9976 ( .C (clk), .D (new_AGEMA_signal_22699), .Q (new_AGEMA_signal_22700) ) ;
    buf_clk new_AGEMA_reg_buffer_9980 ( .C (clk), .D (new_AGEMA_signal_22703), .Q (new_AGEMA_signal_22704) ) ;
    buf_clk new_AGEMA_reg_buffer_9984 ( .C (clk), .D (new_AGEMA_signal_22707), .Q (new_AGEMA_signal_22708) ) ;
    buf_clk new_AGEMA_reg_buffer_9988 ( .C (clk), .D (new_AGEMA_signal_22711), .Q (new_AGEMA_signal_22712) ) ;
    buf_clk new_AGEMA_reg_buffer_9992 ( .C (clk), .D (new_AGEMA_signal_22715), .Q (new_AGEMA_signal_22716) ) ;
    buf_clk new_AGEMA_reg_buffer_9996 ( .C (clk), .D (new_AGEMA_signal_22719), .Q (new_AGEMA_signal_22720) ) ;
    buf_clk new_AGEMA_reg_buffer_10000 ( .C (clk), .D (new_AGEMA_signal_22723), .Q (new_AGEMA_signal_22724) ) ;
    buf_clk new_AGEMA_reg_buffer_10004 ( .C (clk), .D (new_AGEMA_signal_22727), .Q (new_AGEMA_signal_22728) ) ;
    buf_clk new_AGEMA_reg_buffer_10008 ( .C (clk), .D (new_AGEMA_signal_22731), .Q (new_AGEMA_signal_22732) ) ;
    buf_clk new_AGEMA_reg_buffer_10012 ( .C (clk), .D (new_AGEMA_signal_22735), .Q (new_AGEMA_signal_22736) ) ;
    buf_clk new_AGEMA_reg_buffer_10016 ( .C (clk), .D (new_AGEMA_signal_22739), .Q (new_AGEMA_signal_22740) ) ;
    buf_clk new_AGEMA_reg_buffer_10020 ( .C (clk), .D (new_AGEMA_signal_22743), .Q (new_AGEMA_signal_22744) ) ;
    buf_clk new_AGEMA_reg_buffer_10024 ( .C (clk), .D (new_AGEMA_signal_22747), .Q (new_AGEMA_signal_22748) ) ;
    buf_clk new_AGEMA_reg_buffer_10028 ( .C (clk), .D (new_AGEMA_signal_22751), .Q (new_AGEMA_signal_22752) ) ;
    buf_clk new_AGEMA_reg_buffer_10032 ( .C (clk), .D (new_AGEMA_signal_22755), .Q (new_AGEMA_signal_22756) ) ;
    buf_clk new_AGEMA_reg_buffer_10036 ( .C (clk), .D (new_AGEMA_signal_22759), .Q (new_AGEMA_signal_22760) ) ;
    buf_clk new_AGEMA_reg_buffer_10040 ( .C (clk), .D (new_AGEMA_signal_22763), .Q (new_AGEMA_signal_22764) ) ;
    buf_clk new_AGEMA_reg_buffer_10044 ( .C (clk), .D (new_AGEMA_signal_22767), .Q (new_AGEMA_signal_22768) ) ;
    buf_clk new_AGEMA_reg_buffer_10048 ( .C (clk), .D (new_AGEMA_signal_22771), .Q (new_AGEMA_signal_22772) ) ;
    buf_clk new_AGEMA_reg_buffer_10052 ( .C (clk), .D (new_AGEMA_signal_22775), .Q (new_AGEMA_signal_22776) ) ;
    buf_clk new_AGEMA_reg_buffer_10056 ( .C (clk), .D (new_AGEMA_signal_22779), .Q (new_AGEMA_signal_22780) ) ;
    buf_clk new_AGEMA_reg_buffer_10060 ( .C (clk), .D (new_AGEMA_signal_22783), .Q (new_AGEMA_signal_22784) ) ;
    buf_clk new_AGEMA_reg_buffer_10064 ( .C (clk), .D (new_AGEMA_signal_22787), .Q (new_AGEMA_signal_22788) ) ;
    buf_clk new_AGEMA_reg_buffer_10068 ( .C (clk), .D (new_AGEMA_signal_22791), .Q (new_AGEMA_signal_22792) ) ;
    buf_clk new_AGEMA_reg_buffer_10072 ( .C (clk), .D (new_AGEMA_signal_22795), .Q (new_AGEMA_signal_22796) ) ;
    buf_clk new_AGEMA_reg_buffer_10076 ( .C (clk), .D (new_AGEMA_signal_22799), .Q (new_AGEMA_signal_22800) ) ;
    buf_clk new_AGEMA_reg_buffer_10080 ( .C (clk), .D (new_AGEMA_signal_22803), .Q (new_AGEMA_signal_22804) ) ;
    buf_clk new_AGEMA_reg_buffer_10084 ( .C (clk), .D (new_AGEMA_signal_22807), .Q (new_AGEMA_signal_22808) ) ;
    buf_clk new_AGEMA_reg_buffer_10088 ( .C (clk), .D (new_AGEMA_signal_22811), .Q (new_AGEMA_signal_22812) ) ;
    buf_clk new_AGEMA_reg_buffer_10092 ( .C (clk), .D (new_AGEMA_signal_22815), .Q (new_AGEMA_signal_22816) ) ;
    buf_clk new_AGEMA_reg_buffer_10096 ( .C (clk), .D (new_AGEMA_signal_22819), .Q (new_AGEMA_signal_22820) ) ;
    buf_clk new_AGEMA_reg_buffer_10100 ( .C (clk), .D (new_AGEMA_signal_22823), .Q (new_AGEMA_signal_22824) ) ;
    buf_clk new_AGEMA_reg_buffer_10104 ( .C (clk), .D (new_AGEMA_signal_22827), .Q (new_AGEMA_signal_22828) ) ;
    buf_clk new_AGEMA_reg_buffer_10108 ( .C (clk), .D (new_AGEMA_signal_22831), .Q (new_AGEMA_signal_22832) ) ;
    buf_clk new_AGEMA_reg_buffer_10112 ( .C (clk), .D (new_AGEMA_signal_22835), .Q (new_AGEMA_signal_22836) ) ;
    buf_clk new_AGEMA_reg_buffer_10116 ( .C (clk), .D (new_AGEMA_signal_22839), .Q (new_AGEMA_signal_22840) ) ;
    buf_clk new_AGEMA_reg_buffer_10120 ( .C (clk), .D (new_AGEMA_signal_22843), .Q (new_AGEMA_signal_22844) ) ;
    buf_clk new_AGEMA_reg_buffer_10124 ( .C (clk), .D (new_AGEMA_signal_22847), .Q (new_AGEMA_signal_22848) ) ;
    buf_clk new_AGEMA_reg_buffer_10128 ( .C (clk), .D (new_AGEMA_signal_22851), .Q (new_AGEMA_signal_22852) ) ;
    buf_clk new_AGEMA_reg_buffer_10132 ( .C (clk), .D (new_AGEMA_signal_22855), .Q (new_AGEMA_signal_22856) ) ;
    buf_clk new_AGEMA_reg_buffer_10136 ( .C (clk), .D (new_AGEMA_signal_22859), .Q (new_AGEMA_signal_22860) ) ;
    buf_clk new_AGEMA_reg_buffer_10140 ( .C (clk), .D (new_AGEMA_signal_22863), .Q (new_AGEMA_signal_22864) ) ;
    buf_clk new_AGEMA_reg_buffer_10144 ( .C (clk), .D (new_AGEMA_signal_22867), .Q (new_AGEMA_signal_22868) ) ;
    buf_clk new_AGEMA_reg_buffer_10148 ( .C (clk), .D (new_AGEMA_signal_22871), .Q (new_AGEMA_signal_22872) ) ;
    buf_clk new_AGEMA_reg_buffer_10152 ( .C (clk), .D (new_AGEMA_signal_22875), .Q (new_AGEMA_signal_22876) ) ;
    buf_clk new_AGEMA_reg_buffer_10156 ( .C (clk), .D (new_AGEMA_signal_22879), .Q (new_AGEMA_signal_22880) ) ;
    buf_clk new_AGEMA_reg_buffer_10160 ( .C (clk), .D (new_AGEMA_signal_22883), .Q (new_AGEMA_signal_22884) ) ;
    buf_clk new_AGEMA_reg_buffer_10164 ( .C (clk), .D (new_AGEMA_signal_22887), .Q (new_AGEMA_signal_22888) ) ;
    buf_clk new_AGEMA_reg_buffer_10168 ( .C (clk), .D (new_AGEMA_signal_22891), .Q (new_AGEMA_signal_22892) ) ;
    buf_clk new_AGEMA_reg_buffer_10172 ( .C (clk), .D (new_AGEMA_signal_22895), .Q (new_AGEMA_signal_22896) ) ;
    buf_clk new_AGEMA_reg_buffer_10176 ( .C (clk), .D (new_AGEMA_signal_22899), .Q (new_AGEMA_signal_22900) ) ;
    buf_clk new_AGEMA_reg_buffer_10180 ( .C (clk), .D (new_AGEMA_signal_22903), .Q (new_AGEMA_signal_22904) ) ;
    buf_clk new_AGEMA_reg_buffer_10184 ( .C (clk), .D (new_AGEMA_signal_22907), .Q (new_AGEMA_signal_22908) ) ;
    buf_clk new_AGEMA_reg_buffer_10188 ( .C (clk), .D (new_AGEMA_signal_22911), .Q (new_AGEMA_signal_22912) ) ;
    buf_clk new_AGEMA_reg_buffer_10192 ( .C (clk), .D (new_AGEMA_signal_22915), .Q (new_AGEMA_signal_22916) ) ;
    buf_clk new_AGEMA_reg_buffer_10196 ( .C (clk), .D (new_AGEMA_signal_22919), .Q (new_AGEMA_signal_22920) ) ;
    buf_clk new_AGEMA_reg_buffer_10200 ( .C (clk), .D (new_AGEMA_signal_22923), .Q (new_AGEMA_signal_22924) ) ;
    buf_clk new_AGEMA_reg_buffer_10204 ( .C (clk), .D (new_AGEMA_signal_22927), .Q (new_AGEMA_signal_22928) ) ;
    buf_clk new_AGEMA_reg_buffer_10208 ( .C (clk), .D (new_AGEMA_signal_22931), .Q (new_AGEMA_signal_22932) ) ;
    buf_clk new_AGEMA_reg_buffer_10212 ( .C (clk), .D (new_AGEMA_signal_22935), .Q (new_AGEMA_signal_22936) ) ;
    buf_clk new_AGEMA_reg_buffer_10216 ( .C (clk), .D (new_AGEMA_signal_22939), .Q (new_AGEMA_signal_22940) ) ;
    buf_clk new_AGEMA_reg_buffer_10220 ( .C (clk), .D (new_AGEMA_signal_22943), .Q (new_AGEMA_signal_22944) ) ;
    buf_clk new_AGEMA_reg_buffer_10224 ( .C (clk), .D (new_AGEMA_signal_22947), .Q (new_AGEMA_signal_22948) ) ;
    buf_clk new_AGEMA_reg_buffer_10228 ( .C (clk), .D (new_AGEMA_signal_22951), .Q (new_AGEMA_signal_22952) ) ;
    buf_clk new_AGEMA_reg_buffer_10232 ( .C (clk), .D (new_AGEMA_signal_22955), .Q (new_AGEMA_signal_22956) ) ;
    buf_clk new_AGEMA_reg_buffer_10236 ( .C (clk), .D (new_AGEMA_signal_22959), .Q (new_AGEMA_signal_22960) ) ;
    buf_clk new_AGEMA_reg_buffer_10240 ( .C (clk), .D (new_AGEMA_signal_22963), .Q (new_AGEMA_signal_22964) ) ;
    buf_clk new_AGEMA_reg_buffer_10244 ( .C (clk), .D (new_AGEMA_signal_22967), .Q (new_AGEMA_signal_22968) ) ;
    buf_clk new_AGEMA_reg_buffer_10248 ( .C (clk), .D (new_AGEMA_signal_22971), .Q (new_AGEMA_signal_22972) ) ;
    buf_clk new_AGEMA_reg_buffer_10252 ( .C (clk), .D (new_AGEMA_signal_22975), .Q (new_AGEMA_signal_22976) ) ;
    buf_clk new_AGEMA_reg_buffer_10256 ( .C (clk), .D (new_AGEMA_signal_22979), .Q (new_AGEMA_signal_22980) ) ;
    buf_clk new_AGEMA_reg_buffer_10260 ( .C (clk), .D (new_AGEMA_signal_22983), .Q (new_AGEMA_signal_22984) ) ;
    buf_clk new_AGEMA_reg_buffer_10264 ( .C (clk), .D (new_AGEMA_signal_22987), .Q (new_AGEMA_signal_22988) ) ;
    buf_clk new_AGEMA_reg_buffer_10268 ( .C (clk), .D (new_AGEMA_signal_22991), .Q (new_AGEMA_signal_22992) ) ;
    buf_clk new_AGEMA_reg_buffer_10272 ( .C (clk), .D (new_AGEMA_signal_22995), .Q (new_AGEMA_signal_22996) ) ;
    buf_clk new_AGEMA_reg_buffer_10276 ( .C (clk), .D (new_AGEMA_signal_22999), .Q (new_AGEMA_signal_23000) ) ;
    buf_clk new_AGEMA_reg_buffer_10280 ( .C (clk), .D (new_AGEMA_signal_23003), .Q (new_AGEMA_signal_23004) ) ;
    buf_clk new_AGEMA_reg_buffer_10284 ( .C (clk), .D (new_AGEMA_signal_23007), .Q (new_AGEMA_signal_23008) ) ;
    buf_clk new_AGEMA_reg_buffer_10288 ( .C (clk), .D (new_AGEMA_signal_23011), .Q (new_AGEMA_signal_23012) ) ;
    buf_clk new_AGEMA_reg_buffer_10292 ( .C (clk), .D (new_AGEMA_signal_23015), .Q (new_AGEMA_signal_23016) ) ;
    buf_clk new_AGEMA_reg_buffer_10296 ( .C (clk), .D (new_AGEMA_signal_23019), .Q (new_AGEMA_signal_23020) ) ;
    buf_clk new_AGEMA_reg_buffer_10300 ( .C (clk), .D (new_AGEMA_signal_23023), .Q (new_AGEMA_signal_23024) ) ;
    buf_clk new_AGEMA_reg_buffer_10304 ( .C (clk), .D (new_AGEMA_signal_23027), .Q (new_AGEMA_signal_23028) ) ;
    buf_clk new_AGEMA_reg_buffer_10308 ( .C (clk), .D (new_AGEMA_signal_23031), .Q (new_AGEMA_signal_23032) ) ;
    buf_clk new_AGEMA_reg_buffer_10312 ( .C (clk), .D (new_AGEMA_signal_23035), .Q (new_AGEMA_signal_23036) ) ;
    buf_clk new_AGEMA_reg_buffer_10316 ( .C (clk), .D (new_AGEMA_signal_23039), .Q (new_AGEMA_signal_23040) ) ;
    buf_clk new_AGEMA_reg_buffer_10320 ( .C (clk), .D (new_AGEMA_signal_23043), .Q (new_AGEMA_signal_23044) ) ;
    buf_clk new_AGEMA_reg_buffer_10324 ( .C (clk), .D (new_AGEMA_signal_23047), .Q (new_AGEMA_signal_23048) ) ;
    buf_clk new_AGEMA_reg_buffer_10328 ( .C (clk), .D (new_AGEMA_signal_23051), .Q (new_AGEMA_signal_23052) ) ;
    buf_clk new_AGEMA_reg_buffer_10332 ( .C (clk), .D (new_AGEMA_signal_23055), .Q (new_AGEMA_signal_23056) ) ;
    buf_clk new_AGEMA_reg_buffer_10336 ( .C (clk), .D (new_AGEMA_signal_23059), .Q (new_AGEMA_signal_23060) ) ;
    buf_clk new_AGEMA_reg_buffer_10340 ( .C (clk), .D (new_AGEMA_signal_23063), .Q (new_AGEMA_signal_23064) ) ;
    buf_clk new_AGEMA_reg_buffer_10344 ( .C (clk), .D (new_AGEMA_signal_23067), .Q (new_AGEMA_signal_23068) ) ;
    buf_clk new_AGEMA_reg_buffer_10348 ( .C (clk), .D (new_AGEMA_signal_23071), .Q (new_AGEMA_signal_23072) ) ;
    buf_clk new_AGEMA_reg_buffer_10352 ( .C (clk), .D (new_AGEMA_signal_23075), .Q (new_AGEMA_signal_23076) ) ;
    buf_clk new_AGEMA_reg_buffer_10356 ( .C (clk), .D (new_AGEMA_signal_23079), .Q (new_AGEMA_signal_23080) ) ;
    buf_clk new_AGEMA_reg_buffer_10360 ( .C (clk), .D (new_AGEMA_signal_23083), .Q (new_AGEMA_signal_23084) ) ;
    buf_clk new_AGEMA_reg_buffer_10364 ( .C (clk), .D (new_AGEMA_signal_23087), .Q (new_AGEMA_signal_23088) ) ;
    buf_clk new_AGEMA_reg_buffer_10368 ( .C (clk), .D (new_AGEMA_signal_23091), .Q (new_AGEMA_signal_23092) ) ;
    buf_clk new_AGEMA_reg_buffer_10372 ( .C (clk), .D (new_AGEMA_signal_23095), .Q (new_AGEMA_signal_23096) ) ;
    buf_clk new_AGEMA_reg_buffer_10376 ( .C (clk), .D (new_AGEMA_signal_23099), .Q (new_AGEMA_signal_23100) ) ;
    buf_clk new_AGEMA_reg_buffer_10380 ( .C (clk), .D (new_AGEMA_signal_23103), .Q (new_AGEMA_signal_23104) ) ;
    buf_clk new_AGEMA_reg_buffer_10384 ( .C (clk), .D (new_AGEMA_signal_23107), .Q (new_AGEMA_signal_23108) ) ;
    buf_clk new_AGEMA_reg_buffer_10388 ( .C (clk), .D (new_AGEMA_signal_23111), .Q (new_AGEMA_signal_23112) ) ;
    buf_clk new_AGEMA_reg_buffer_10392 ( .C (clk), .D (new_AGEMA_signal_23115), .Q (new_AGEMA_signal_23116) ) ;
    buf_clk new_AGEMA_reg_buffer_10396 ( .C (clk), .D (new_AGEMA_signal_23119), .Q (new_AGEMA_signal_23120) ) ;
    buf_clk new_AGEMA_reg_buffer_10400 ( .C (clk), .D (new_AGEMA_signal_23123), .Q (new_AGEMA_signal_23124) ) ;
    buf_clk new_AGEMA_reg_buffer_10404 ( .C (clk), .D (new_AGEMA_signal_23127), .Q (new_AGEMA_signal_23128) ) ;
    buf_clk new_AGEMA_reg_buffer_10408 ( .C (clk), .D (new_AGEMA_signal_23131), .Q (new_AGEMA_signal_23132) ) ;
    buf_clk new_AGEMA_reg_buffer_10412 ( .C (clk), .D (new_AGEMA_signal_23135), .Q (new_AGEMA_signal_23136) ) ;
    buf_clk new_AGEMA_reg_buffer_10416 ( .C (clk), .D (new_AGEMA_signal_23139), .Q (new_AGEMA_signal_23140) ) ;
    buf_clk new_AGEMA_reg_buffer_10420 ( .C (clk), .D (new_AGEMA_signal_23143), .Q (new_AGEMA_signal_23144) ) ;
    buf_clk new_AGEMA_reg_buffer_10424 ( .C (clk), .D (new_AGEMA_signal_23147), .Q (new_AGEMA_signal_23148) ) ;
    buf_clk new_AGEMA_reg_buffer_10428 ( .C (clk), .D (new_AGEMA_signal_23151), .Q (new_AGEMA_signal_23152) ) ;
    buf_clk new_AGEMA_reg_buffer_10432 ( .C (clk), .D (new_AGEMA_signal_23155), .Q (new_AGEMA_signal_23156) ) ;
    buf_clk new_AGEMA_reg_buffer_10436 ( .C (clk), .D (new_AGEMA_signal_23159), .Q (new_AGEMA_signal_23160) ) ;
    buf_clk new_AGEMA_reg_buffer_10440 ( .C (clk), .D (new_AGEMA_signal_23163), .Q (new_AGEMA_signal_23164) ) ;
    buf_clk new_AGEMA_reg_buffer_10444 ( .C (clk), .D (new_AGEMA_signal_23167), .Q (new_AGEMA_signal_23168) ) ;
    buf_clk new_AGEMA_reg_buffer_10448 ( .C (clk), .D (new_AGEMA_signal_23171), .Q (new_AGEMA_signal_23172) ) ;
    buf_clk new_AGEMA_reg_buffer_10452 ( .C (clk), .D (new_AGEMA_signal_23175), .Q (new_AGEMA_signal_23176) ) ;
    buf_clk new_AGEMA_reg_buffer_10456 ( .C (clk), .D (new_AGEMA_signal_23179), .Q (new_AGEMA_signal_23180) ) ;
    buf_clk new_AGEMA_reg_buffer_10460 ( .C (clk), .D (new_AGEMA_signal_23183), .Q (new_AGEMA_signal_23184) ) ;
    buf_clk new_AGEMA_reg_buffer_10464 ( .C (clk), .D (new_AGEMA_signal_23187), .Q (new_AGEMA_signal_23188) ) ;
    buf_clk new_AGEMA_reg_buffer_10468 ( .C (clk), .D (new_AGEMA_signal_23191), .Q (new_AGEMA_signal_23192) ) ;
    buf_clk new_AGEMA_reg_buffer_10472 ( .C (clk), .D (new_AGEMA_signal_23195), .Q (new_AGEMA_signal_23196) ) ;
    buf_clk new_AGEMA_reg_buffer_10476 ( .C (clk), .D (new_AGEMA_signal_23199), .Q (new_AGEMA_signal_23200) ) ;
    buf_clk new_AGEMA_reg_buffer_10480 ( .C (clk), .D (new_AGEMA_signal_23203), .Q (new_AGEMA_signal_23204) ) ;
    buf_clk new_AGEMA_reg_buffer_10484 ( .C (clk), .D (new_AGEMA_signal_23207), .Q (new_AGEMA_signal_23208) ) ;
    buf_clk new_AGEMA_reg_buffer_10488 ( .C (clk), .D (new_AGEMA_signal_23211), .Q (new_AGEMA_signal_23212) ) ;
    buf_clk new_AGEMA_reg_buffer_10492 ( .C (clk), .D (new_AGEMA_signal_23215), .Q (new_AGEMA_signal_23216) ) ;
    buf_clk new_AGEMA_reg_buffer_10496 ( .C (clk), .D (new_AGEMA_signal_23219), .Q (new_AGEMA_signal_23220) ) ;
    buf_clk new_AGEMA_reg_buffer_10500 ( .C (clk), .D (new_AGEMA_signal_23223), .Q (new_AGEMA_signal_23224) ) ;
    buf_clk new_AGEMA_reg_buffer_10504 ( .C (clk), .D (new_AGEMA_signal_23227), .Q (new_AGEMA_signal_23228) ) ;
    buf_clk new_AGEMA_reg_buffer_10508 ( .C (clk), .D (new_AGEMA_signal_23231), .Q (new_AGEMA_signal_23232) ) ;
    buf_clk new_AGEMA_reg_buffer_10512 ( .C (clk), .D (new_AGEMA_signal_23235), .Q (new_AGEMA_signal_23236) ) ;
    buf_clk new_AGEMA_reg_buffer_10516 ( .C (clk), .D (new_AGEMA_signal_23239), .Q (new_AGEMA_signal_23240) ) ;
    buf_clk new_AGEMA_reg_buffer_10520 ( .C (clk), .D (new_AGEMA_signal_23243), .Q (new_AGEMA_signal_23244) ) ;
    buf_clk new_AGEMA_reg_buffer_10524 ( .C (clk), .D (new_AGEMA_signal_23247), .Q (new_AGEMA_signal_23248) ) ;
    buf_clk new_AGEMA_reg_buffer_10528 ( .C (clk), .D (new_AGEMA_signal_23251), .Q (new_AGEMA_signal_23252) ) ;
    buf_clk new_AGEMA_reg_buffer_10532 ( .C (clk), .D (new_AGEMA_signal_23255), .Q (new_AGEMA_signal_23256) ) ;
    buf_clk new_AGEMA_reg_buffer_10536 ( .C (clk), .D (new_AGEMA_signal_23259), .Q (new_AGEMA_signal_23260) ) ;
    buf_clk new_AGEMA_reg_buffer_10540 ( .C (clk), .D (new_AGEMA_signal_23263), .Q (new_AGEMA_signal_23264) ) ;
    buf_clk new_AGEMA_reg_buffer_10544 ( .C (clk), .D (new_AGEMA_signal_23267), .Q (new_AGEMA_signal_23268) ) ;
    buf_clk new_AGEMA_reg_buffer_10548 ( .C (clk), .D (new_AGEMA_signal_23271), .Q (new_AGEMA_signal_23272) ) ;
    buf_clk new_AGEMA_reg_buffer_10552 ( .C (clk), .D (new_AGEMA_signal_23275), .Q (new_AGEMA_signal_23276) ) ;
    buf_clk new_AGEMA_reg_buffer_10556 ( .C (clk), .D (new_AGEMA_signal_23279), .Q (new_AGEMA_signal_23280) ) ;
    buf_clk new_AGEMA_reg_buffer_10560 ( .C (clk), .D (new_AGEMA_signal_23283), .Q (new_AGEMA_signal_23284) ) ;
    buf_clk new_AGEMA_reg_buffer_10564 ( .C (clk), .D (new_AGEMA_signal_23287), .Q (new_AGEMA_signal_23288) ) ;
    buf_clk new_AGEMA_reg_buffer_10568 ( .C (clk), .D (new_AGEMA_signal_23291), .Q (new_AGEMA_signal_23292) ) ;
    buf_clk new_AGEMA_reg_buffer_10572 ( .C (clk), .D (new_AGEMA_signal_23295), .Q (new_AGEMA_signal_23296) ) ;
    buf_clk new_AGEMA_reg_buffer_10576 ( .C (clk), .D (new_AGEMA_signal_23299), .Q (new_AGEMA_signal_23300) ) ;
    buf_clk new_AGEMA_reg_buffer_10580 ( .C (clk), .D (new_AGEMA_signal_23303), .Q (new_AGEMA_signal_23304) ) ;
    buf_clk new_AGEMA_reg_buffer_10584 ( .C (clk), .D (new_AGEMA_signal_23307), .Q (new_AGEMA_signal_23308) ) ;
    buf_clk new_AGEMA_reg_buffer_10588 ( .C (clk), .D (new_AGEMA_signal_23311), .Q (new_AGEMA_signal_23312) ) ;
    buf_clk new_AGEMA_reg_buffer_10592 ( .C (clk), .D (new_AGEMA_signal_23315), .Q (new_AGEMA_signal_23316) ) ;
    buf_clk new_AGEMA_reg_buffer_10596 ( .C (clk), .D (new_AGEMA_signal_23319), .Q (new_AGEMA_signal_23320) ) ;
    buf_clk new_AGEMA_reg_buffer_10600 ( .C (clk), .D (new_AGEMA_signal_23323), .Q (new_AGEMA_signal_23324) ) ;
    buf_clk new_AGEMA_reg_buffer_10604 ( .C (clk), .D (new_AGEMA_signal_23327), .Q (new_AGEMA_signal_23328) ) ;
    buf_clk new_AGEMA_reg_buffer_10608 ( .C (clk), .D (new_AGEMA_signal_23331), .Q (new_AGEMA_signal_23332) ) ;
    buf_clk new_AGEMA_reg_buffer_10612 ( .C (clk), .D (new_AGEMA_signal_23335), .Q (new_AGEMA_signal_23336) ) ;
    buf_clk new_AGEMA_reg_buffer_10616 ( .C (clk), .D (new_AGEMA_signal_23339), .Q (new_AGEMA_signal_23340) ) ;
    buf_clk new_AGEMA_reg_buffer_10620 ( .C (clk), .D (new_AGEMA_signal_23343), .Q (new_AGEMA_signal_23344) ) ;
    buf_clk new_AGEMA_reg_buffer_10624 ( .C (clk), .D (new_AGEMA_signal_23347), .Q (new_AGEMA_signal_23348) ) ;
    buf_clk new_AGEMA_reg_buffer_10628 ( .C (clk), .D (new_AGEMA_signal_23351), .Q (new_AGEMA_signal_23352) ) ;
    buf_clk new_AGEMA_reg_buffer_10632 ( .C (clk), .D (new_AGEMA_signal_23355), .Q (new_AGEMA_signal_23356) ) ;
    buf_clk new_AGEMA_reg_buffer_10636 ( .C (clk), .D (new_AGEMA_signal_23359), .Q (new_AGEMA_signal_23360) ) ;
    buf_clk new_AGEMA_reg_buffer_10640 ( .C (clk), .D (new_AGEMA_signal_23363), .Q (new_AGEMA_signal_23364) ) ;
    buf_clk new_AGEMA_reg_buffer_10644 ( .C (clk), .D (new_AGEMA_signal_23367), .Q (new_AGEMA_signal_23368) ) ;
    buf_clk new_AGEMA_reg_buffer_10648 ( .C (clk), .D (new_AGEMA_signal_23371), .Q (new_AGEMA_signal_23372) ) ;
    buf_clk new_AGEMA_reg_buffer_10652 ( .C (clk), .D (new_AGEMA_signal_23375), .Q (new_AGEMA_signal_23376) ) ;
    buf_clk new_AGEMA_reg_buffer_10656 ( .C (clk), .D (new_AGEMA_signal_23379), .Q (new_AGEMA_signal_23380) ) ;
    buf_clk new_AGEMA_reg_buffer_10660 ( .C (clk), .D (new_AGEMA_signal_23383), .Q (new_AGEMA_signal_23384) ) ;
    buf_clk new_AGEMA_reg_buffer_10664 ( .C (clk), .D (new_AGEMA_signal_23387), .Q (new_AGEMA_signal_23388) ) ;
    buf_clk new_AGEMA_reg_buffer_10668 ( .C (clk), .D (new_AGEMA_signal_23391), .Q (new_AGEMA_signal_23392) ) ;
    buf_clk new_AGEMA_reg_buffer_10672 ( .C (clk), .D (new_AGEMA_signal_23395), .Q (new_AGEMA_signal_23396) ) ;
    buf_clk new_AGEMA_reg_buffer_10676 ( .C (clk), .D (new_AGEMA_signal_23399), .Q (new_AGEMA_signal_23400) ) ;
    buf_clk new_AGEMA_reg_buffer_10680 ( .C (clk), .D (new_AGEMA_signal_23403), .Q (new_AGEMA_signal_23404) ) ;
    buf_clk new_AGEMA_reg_buffer_10684 ( .C (clk), .D (new_AGEMA_signal_23407), .Q (new_AGEMA_signal_23408) ) ;
    buf_clk new_AGEMA_reg_buffer_10688 ( .C (clk), .D (new_AGEMA_signal_23411), .Q (new_AGEMA_signal_23412) ) ;
    buf_clk new_AGEMA_reg_buffer_10692 ( .C (clk), .D (new_AGEMA_signal_23415), .Q (new_AGEMA_signal_23416) ) ;
    buf_clk new_AGEMA_reg_buffer_10696 ( .C (clk), .D (new_AGEMA_signal_23419), .Q (new_AGEMA_signal_23420) ) ;
    buf_clk new_AGEMA_reg_buffer_10700 ( .C (clk), .D (new_AGEMA_signal_23423), .Q (new_AGEMA_signal_23424) ) ;
    buf_clk new_AGEMA_reg_buffer_10704 ( .C (clk), .D (new_AGEMA_signal_23427), .Q (new_AGEMA_signal_23428) ) ;
    buf_clk new_AGEMA_reg_buffer_10708 ( .C (clk), .D (new_AGEMA_signal_23431), .Q (new_AGEMA_signal_23432) ) ;
    buf_clk new_AGEMA_reg_buffer_10712 ( .C (clk), .D (new_AGEMA_signal_23435), .Q (new_AGEMA_signal_23436) ) ;
    buf_clk new_AGEMA_reg_buffer_10716 ( .C (clk), .D (new_AGEMA_signal_23439), .Q (new_AGEMA_signal_23440) ) ;
    buf_clk new_AGEMA_reg_buffer_10720 ( .C (clk), .D (new_AGEMA_signal_23443), .Q (new_AGEMA_signal_23444) ) ;
    buf_clk new_AGEMA_reg_buffer_10724 ( .C (clk), .D (new_AGEMA_signal_23447), .Q (new_AGEMA_signal_23448) ) ;
    buf_clk new_AGEMA_reg_buffer_10728 ( .C (clk), .D (new_AGEMA_signal_23451), .Q (new_AGEMA_signal_23452) ) ;
    buf_clk new_AGEMA_reg_buffer_10732 ( .C (clk), .D (new_AGEMA_signal_23455), .Q (new_AGEMA_signal_23456) ) ;
    buf_clk new_AGEMA_reg_buffer_10736 ( .C (clk), .D (new_AGEMA_signal_23459), .Q (new_AGEMA_signal_23460) ) ;
    buf_clk new_AGEMA_reg_buffer_10740 ( .C (clk), .D (new_AGEMA_signal_23463), .Q (new_AGEMA_signal_23464) ) ;
    buf_clk new_AGEMA_reg_buffer_10744 ( .C (clk), .D (new_AGEMA_signal_23467), .Q (new_AGEMA_signal_23468) ) ;
    buf_clk new_AGEMA_reg_buffer_10748 ( .C (clk), .D (new_AGEMA_signal_23471), .Q (new_AGEMA_signal_23472) ) ;
    buf_clk new_AGEMA_reg_buffer_10752 ( .C (clk), .D (new_AGEMA_signal_23475), .Q (new_AGEMA_signal_23476) ) ;
    buf_clk new_AGEMA_reg_buffer_10756 ( .C (clk), .D (new_AGEMA_signal_23479), .Q (new_AGEMA_signal_23480) ) ;
    buf_clk new_AGEMA_reg_buffer_10760 ( .C (clk), .D (new_AGEMA_signal_23483), .Q (new_AGEMA_signal_23484) ) ;
    buf_clk new_AGEMA_reg_buffer_10764 ( .C (clk), .D (new_AGEMA_signal_23487), .Q (new_AGEMA_signal_23488) ) ;
    buf_clk new_AGEMA_reg_buffer_10768 ( .C (clk), .D (new_AGEMA_signal_23491), .Q (new_AGEMA_signal_23492) ) ;
    buf_clk new_AGEMA_reg_buffer_10772 ( .C (clk), .D (new_AGEMA_signal_23495), .Q (new_AGEMA_signal_23496) ) ;
    buf_clk new_AGEMA_reg_buffer_10776 ( .C (clk), .D (new_AGEMA_signal_23499), .Q (new_AGEMA_signal_23500) ) ;
    buf_clk new_AGEMA_reg_buffer_10780 ( .C (clk), .D (new_AGEMA_signal_23503), .Q (new_AGEMA_signal_23504) ) ;
    buf_clk new_AGEMA_reg_buffer_10784 ( .C (clk), .D (new_AGEMA_signal_23507), .Q (new_AGEMA_signal_23508) ) ;
    buf_clk new_AGEMA_reg_buffer_10788 ( .C (clk), .D (new_AGEMA_signal_23511), .Q (new_AGEMA_signal_23512) ) ;
    buf_clk new_AGEMA_reg_buffer_10792 ( .C (clk), .D (new_AGEMA_signal_23515), .Q (new_AGEMA_signal_23516) ) ;
    buf_clk new_AGEMA_reg_buffer_10796 ( .C (clk), .D (new_AGEMA_signal_23519), .Q (new_AGEMA_signal_23520) ) ;
    buf_clk new_AGEMA_reg_buffer_10800 ( .C (clk), .D (new_AGEMA_signal_23523), .Q (new_AGEMA_signal_23524) ) ;
    buf_clk new_AGEMA_reg_buffer_10804 ( .C (clk), .D (new_AGEMA_signal_23527), .Q (new_AGEMA_signal_23528) ) ;
    buf_clk new_AGEMA_reg_buffer_10808 ( .C (clk), .D (new_AGEMA_signal_23531), .Q (new_AGEMA_signal_23532) ) ;
    buf_clk new_AGEMA_reg_buffer_10812 ( .C (clk), .D (new_AGEMA_signal_23535), .Q (new_AGEMA_signal_23536) ) ;
    buf_clk new_AGEMA_reg_buffer_10816 ( .C (clk), .D (new_AGEMA_signal_23539), .Q (new_AGEMA_signal_23540) ) ;
    buf_clk new_AGEMA_reg_buffer_10820 ( .C (clk), .D (new_AGEMA_signal_23543), .Q (new_AGEMA_signal_23544) ) ;
    buf_clk new_AGEMA_reg_buffer_10824 ( .C (clk), .D (new_AGEMA_signal_23547), .Q (new_AGEMA_signal_23548) ) ;
    buf_clk new_AGEMA_reg_buffer_10828 ( .C (clk), .D (new_AGEMA_signal_23551), .Q (new_AGEMA_signal_23552) ) ;
    buf_clk new_AGEMA_reg_buffer_10832 ( .C (clk), .D (new_AGEMA_signal_23555), .Q (new_AGEMA_signal_23556) ) ;
    buf_clk new_AGEMA_reg_buffer_10836 ( .C (clk), .D (new_AGEMA_signal_23559), .Q (new_AGEMA_signal_23560) ) ;
    buf_clk new_AGEMA_reg_buffer_10840 ( .C (clk), .D (new_AGEMA_signal_23563), .Q (new_AGEMA_signal_23564) ) ;
    buf_clk new_AGEMA_reg_buffer_10844 ( .C (clk), .D (new_AGEMA_signal_23567), .Q (new_AGEMA_signal_23568) ) ;
    buf_clk new_AGEMA_reg_buffer_10848 ( .C (clk), .D (new_AGEMA_signal_23571), .Q (new_AGEMA_signal_23572) ) ;
    buf_clk new_AGEMA_reg_buffer_10852 ( .C (clk), .D (new_AGEMA_signal_23575), .Q (new_AGEMA_signal_23576) ) ;
    buf_clk new_AGEMA_reg_buffer_10856 ( .C (clk), .D (new_AGEMA_signal_23579), .Q (new_AGEMA_signal_23580) ) ;
    buf_clk new_AGEMA_reg_buffer_10860 ( .C (clk), .D (new_AGEMA_signal_23583), .Q (new_AGEMA_signal_23584) ) ;
    buf_clk new_AGEMA_reg_buffer_10864 ( .C (clk), .D (new_AGEMA_signal_23587), .Q (new_AGEMA_signal_23588) ) ;
    buf_clk new_AGEMA_reg_buffer_10868 ( .C (clk), .D (new_AGEMA_signal_23591), .Q (new_AGEMA_signal_23592) ) ;
    buf_clk new_AGEMA_reg_buffer_10872 ( .C (clk), .D (new_AGEMA_signal_23595), .Q (new_AGEMA_signal_23596) ) ;
    buf_clk new_AGEMA_reg_buffer_10876 ( .C (clk), .D (new_AGEMA_signal_23599), .Q (new_AGEMA_signal_23600) ) ;
    buf_clk new_AGEMA_reg_buffer_10880 ( .C (clk), .D (new_AGEMA_signal_23603), .Q (new_AGEMA_signal_23604) ) ;
    buf_clk new_AGEMA_reg_buffer_10884 ( .C (clk), .D (new_AGEMA_signal_23607), .Q (new_AGEMA_signal_23608) ) ;
    buf_clk new_AGEMA_reg_buffer_10888 ( .C (clk), .D (new_AGEMA_signal_23611), .Q (new_AGEMA_signal_23612) ) ;
    buf_clk new_AGEMA_reg_buffer_10892 ( .C (clk), .D (new_AGEMA_signal_23615), .Q (new_AGEMA_signal_23616) ) ;
    buf_clk new_AGEMA_reg_buffer_10896 ( .C (clk), .D (new_AGEMA_signal_23619), .Q (new_AGEMA_signal_23620) ) ;
    buf_clk new_AGEMA_reg_buffer_10900 ( .C (clk), .D (new_AGEMA_signal_23623), .Q (new_AGEMA_signal_23624) ) ;
    buf_clk new_AGEMA_reg_buffer_10904 ( .C (clk), .D (new_AGEMA_signal_23627), .Q (new_AGEMA_signal_23628) ) ;
    buf_clk new_AGEMA_reg_buffer_10908 ( .C (clk), .D (new_AGEMA_signal_23631), .Q (new_AGEMA_signal_23632) ) ;
    buf_clk new_AGEMA_reg_buffer_10912 ( .C (clk), .D (new_AGEMA_signal_23635), .Q (new_AGEMA_signal_23636) ) ;
    buf_clk new_AGEMA_reg_buffer_10916 ( .C (clk), .D (new_AGEMA_signal_23639), .Q (new_AGEMA_signal_23640) ) ;
    buf_clk new_AGEMA_reg_buffer_10920 ( .C (clk), .D (new_AGEMA_signal_23643), .Q (new_AGEMA_signal_23644) ) ;
    buf_clk new_AGEMA_reg_buffer_10924 ( .C (clk), .D (new_AGEMA_signal_23647), .Q (new_AGEMA_signal_23648) ) ;
    buf_clk new_AGEMA_reg_buffer_10928 ( .C (clk), .D (new_AGEMA_signal_23651), .Q (new_AGEMA_signal_23652) ) ;
    buf_clk new_AGEMA_reg_buffer_10932 ( .C (clk), .D (new_AGEMA_signal_23655), .Q (new_AGEMA_signal_23656) ) ;
    buf_clk new_AGEMA_reg_buffer_10936 ( .C (clk), .D (new_AGEMA_signal_23659), .Q (new_AGEMA_signal_23660) ) ;
    buf_clk new_AGEMA_reg_buffer_10940 ( .C (clk), .D (new_AGEMA_signal_23663), .Q (new_AGEMA_signal_23664) ) ;
    buf_clk new_AGEMA_reg_buffer_10944 ( .C (clk), .D (new_AGEMA_signal_23667), .Q (new_AGEMA_signal_23668) ) ;
    buf_clk new_AGEMA_reg_buffer_10948 ( .C (clk), .D (new_AGEMA_signal_23671), .Q (new_AGEMA_signal_23672) ) ;
    buf_clk new_AGEMA_reg_buffer_10952 ( .C (clk), .D (new_AGEMA_signal_23675), .Q (new_AGEMA_signal_23676) ) ;
    buf_clk new_AGEMA_reg_buffer_10956 ( .C (clk), .D (new_AGEMA_signal_23679), .Q (new_AGEMA_signal_23680) ) ;
    buf_clk new_AGEMA_reg_buffer_10960 ( .C (clk), .D (new_AGEMA_signal_23683), .Q (new_AGEMA_signal_23684) ) ;
    buf_clk new_AGEMA_reg_buffer_10964 ( .C (clk), .D (new_AGEMA_signal_23687), .Q (new_AGEMA_signal_23688) ) ;
    buf_clk new_AGEMA_reg_buffer_10968 ( .C (clk), .D (new_AGEMA_signal_23691), .Q (new_AGEMA_signal_23692) ) ;
    buf_clk new_AGEMA_reg_buffer_10972 ( .C (clk), .D (new_AGEMA_signal_23695), .Q (new_AGEMA_signal_23696) ) ;
    buf_clk new_AGEMA_reg_buffer_10976 ( .C (clk), .D (new_AGEMA_signal_23699), .Q (new_AGEMA_signal_23700) ) ;
    buf_clk new_AGEMA_reg_buffer_10980 ( .C (clk), .D (new_AGEMA_signal_23703), .Q (new_AGEMA_signal_23704) ) ;
    buf_clk new_AGEMA_reg_buffer_10984 ( .C (clk), .D (new_AGEMA_signal_23707), .Q (new_AGEMA_signal_23708) ) ;
    buf_clk new_AGEMA_reg_buffer_10988 ( .C (clk), .D (new_AGEMA_signal_23711), .Q (new_AGEMA_signal_23712) ) ;
    buf_clk new_AGEMA_reg_buffer_10992 ( .C (clk), .D (new_AGEMA_signal_23715), .Q (new_AGEMA_signal_23716) ) ;
    buf_clk new_AGEMA_reg_buffer_10996 ( .C (clk), .D (new_AGEMA_signal_23719), .Q (new_AGEMA_signal_23720) ) ;
    buf_clk new_AGEMA_reg_buffer_11000 ( .C (clk), .D (new_AGEMA_signal_23723), .Q (new_AGEMA_signal_23724) ) ;
    buf_clk new_AGEMA_reg_buffer_11004 ( .C (clk), .D (new_AGEMA_signal_23727), .Q (new_AGEMA_signal_23728) ) ;
    buf_clk new_AGEMA_reg_buffer_11008 ( .C (clk), .D (new_AGEMA_signal_23731), .Q (new_AGEMA_signal_23732) ) ;
    buf_clk new_AGEMA_reg_buffer_11012 ( .C (clk), .D (new_AGEMA_signal_23735), .Q (new_AGEMA_signal_23736) ) ;
    buf_clk new_AGEMA_reg_buffer_11016 ( .C (clk), .D (new_AGEMA_signal_23739), .Q (new_AGEMA_signal_23740) ) ;
    buf_clk new_AGEMA_reg_buffer_11020 ( .C (clk), .D (new_AGEMA_signal_23743), .Q (new_AGEMA_signal_23744) ) ;
    buf_clk new_AGEMA_reg_buffer_11024 ( .C (clk), .D (new_AGEMA_signal_23747), .Q (new_AGEMA_signal_23748) ) ;
    buf_clk new_AGEMA_reg_buffer_11028 ( .C (clk), .D (new_AGEMA_signal_23751), .Q (new_AGEMA_signal_23752) ) ;
    buf_clk new_AGEMA_reg_buffer_11032 ( .C (clk), .D (new_AGEMA_signal_23755), .Q (new_AGEMA_signal_23756) ) ;
    buf_clk new_AGEMA_reg_buffer_11036 ( .C (clk), .D (new_AGEMA_signal_23759), .Q (new_AGEMA_signal_23760) ) ;
    buf_clk new_AGEMA_reg_buffer_11040 ( .C (clk), .D (new_AGEMA_signal_23763), .Q (new_AGEMA_signal_23764) ) ;
    buf_clk new_AGEMA_reg_buffer_11044 ( .C (clk), .D (new_AGEMA_signal_23767), .Q (new_AGEMA_signal_23768) ) ;
    buf_clk new_AGEMA_reg_buffer_11048 ( .C (clk), .D (new_AGEMA_signal_23771), .Q (new_AGEMA_signal_23772) ) ;
    buf_clk new_AGEMA_reg_buffer_11052 ( .C (clk), .D (new_AGEMA_signal_23775), .Q (new_AGEMA_signal_23776) ) ;
    buf_clk new_AGEMA_reg_buffer_11056 ( .C (clk), .D (new_AGEMA_signal_23779), .Q (new_AGEMA_signal_23780) ) ;
    buf_clk new_AGEMA_reg_buffer_11060 ( .C (clk), .D (new_AGEMA_signal_23783), .Q (new_AGEMA_signal_23784) ) ;
    buf_clk new_AGEMA_reg_buffer_11064 ( .C (clk), .D (new_AGEMA_signal_23787), .Q (new_AGEMA_signal_23788) ) ;
    buf_clk new_AGEMA_reg_buffer_11068 ( .C (clk), .D (new_AGEMA_signal_23791), .Q (new_AGEMA_signal_23792) ) ;
    buf_clk new_AGEMA_reg_buffer_11072 ( .C (clk), .D (new_AGEMA_signal_23795), .Q (new_AGEMA_signal_23796) ) ;
    buf_clk new_AGEMA_reg_buffer_11076 ( .C (clk), .D (new_AGEMA_signal_23799), .Q (new_AGEMA_signal_23800) ) ;
    buf_clk new_AGEMA_reg_buffer_11080 ( .C (clk), .D (new_AGEMA_signal_23803), .Q (new_AGEMA_signal_23804) ) ;
    buf_clk new_AGEMA_reg_buffer_11084 ( .C (clk), .D (new_AGEMA_signal_23807), .Q (new_AGEMA_signal_23808) ) ;
    buf_clk new_AGEMA_reg_buffer_11088 ( .C (clk), .D (new_AGEMA_signal_23811), .Q (new_AGEMA_signal_23812) ) ;
    buf_clk new_AGEMA_reg_buffer_11092 ( .C (clk), .D (new_AGEMA_signal_23815), .Q (new_AGEMA_signal_23816) ) ;
    buf_clk new_AGEMA_reg_buffer_11096 ( .C (clk), .D (new_AGEMA_signal_23819), .Q (new_AGEMA_signal_23820) ) ;
    buf_clk new_AGEMA_reg_buffer_11100 ( .C (clk), .D (new_AGEMA_signal_23823), .Q (new_AGEMA_signal_23824) ) ;
    buf_clk new_AGEMA_reg_buffer_11104 ( .C (clk), .D (new_AGEMA_signal_23827), .Q (new_AGEMA_signal_23828) ) ;
    buf_clk new_AGEMA_reg_buffer_11108 ( .C (clk), .D (new_AGEMA_signal_23831), .Q (new_AGEMA_signal_23832) ) ;
    buf_clk new_AGEMA_reg_buffer_11112 ( .C (clk), .D (new_AGEMA_signal_23835), .Q (new_AGEMA_signal_23836) ) ;
    buf_clk new_AGEMA_reg_buffer_11116 ( .C (clk), .D (new_AGEMA_signal_23839), .Q (new_AGEMA_signal_23840) ) ;
    buf_clk new_AGEMA_reg_buffer_11120 ( .C (clk), .D (new_AGEMA_signal_23843), .Q (new_AGEMA_signal_23844) ) ;
    buf_clk new_AGEMA_reg_buffer_11124 ( .C (clk), .D (new_AGEMA_signal_23847), .Q (new_AGEMA_signal_23848) ) ;
    buf_clk new_AGEMA_reg_buffer_11128 ( .C (clk), .D (new_AGEMA_signal_23851), .Q (new_AGEMA_signal_23852) ) ;
    buf_clk new_AGEMA_reg_buffer_11132 ( .C (clk), .D (new_AGEMA_signal_23855), .Q (new_AGEMA_signal_23856) ) ;
    buf_clk new_AGEMA_reg_buffer_11136 ( .C (clk), .D (new_AGEMA_signal_23859), .Q (new_AGEMA_signal_23860) ) ;
    buf_clk new_AGEMA_reg_buffer_11140 ( .C (clk), .D (new_AGEMA_signal_23863), .Q (new_AGEMA_signal_23864) ) ;
    buf_clk new_AGEMA_reg_buffer_11144 ( .C (clk), .D (new_AGEMA_signal_23867), .Q (new_AGEMA_signal_23868) ) ;
    buf_clk new_AGEMA_reg_buffer_11148 ( .C (clk), .D (new_AGEMA_signal_23871), .Q (new_AGEMA_signal_23872) ) ;
    buf_clk new_AGEMA_reg_buffer_11152 ( .C (clk), .D (new_AGEMA_signal_23875), .Q (new_AGEMA_signal_23876) ) ;
    buf_clk new_AGEMA_reg_buffer_11156 ( .C (clk), .D (new_AGEMA_signal_23879), .Q (new_AGEMA_signal_23880) ) ;
    buf_clk new_AGEMA_reg_buffer_11160 ( .C (clk), .D (new_AGEMA_signal_23883), .Q (new_AGEMA_signal_23884) ) ;
    buf_clk new_AGEMA_reg_buffer_11164 ( .C (clk), .D (new_AGEMA_signal_23887), .Q (new_AGEMA_signal_23888) ) ;
    buf_clk new_AGEMA_reg_buffer_11168 ( .C (clk), .D (new_AGEMA_signal_23891), .Q (new_AGEMA_signal_23892) ) ;
    buf_clk new_AGEMA_reg_buffer_11172 ( .C (clk), .D (new_AGEMA_signal_23895), .Q (new_AGEMA_signal_23896) ) ;
    buf_clk new_AGEMA_reg_buffer_11176 ( .C (clk), .D (new_AGEMA_signal_23899), .Q (new_AGEMA_signal_23900) ) ;
    buf_clk new_AGEMA_reg_buffer_11180 ( .C (clk), .D (new_AGEMA_signal_23903), .Q (new_AGEMA_signal_23904) ) ;
    buf_clk new_AGEMA_reg_buffer_11184 ( .C (clk), .D (new_AGEMA_signal_23907), .Q (new_AGEMA_signal_23908) ) ;
    buf_clk new_AGEMA_reg_buffer_11188 ( .C (clk), .D (new_AGEMA_signal_23911), .Q (new_AGEMA_signal_23912) ) ;
    buf_clk new_AGEMA_reg_buffer_11192 ( .C (clk), .D (new_AGEMA_signal_23915), .Q (new_AGEMA_signal_23916) ) ;
    buf_clk new_AGEMA_reg_buffer_11196 ( .C (clk), .D (new_AGEMA_signal_23919), .Q (new_AGEMA_signal_23920) ) ;
    buf_clk new_AGEMA_reg_buffer_11200 ( .C (clk), .D (new_AGEMA_signal_23923), .Q (new_AGEMA_signal_23924) ) ;
    buf_clk new_AGEMA_reg_buffer_11204 ( .C (clk), .D (new_AGEMA_signal_23927), .Q (new_AGEMA_signal_23928) ) ;
    buf_clk new_AGEMA_reg_buffer_11208 ( .C (clk), .D (new_AGEMA_signal_23931), .Q (new_AGEMA_signal_23932) ) ;
    buf_clk new_AGEMA_reg_buffer_11212 ( .C (clk), .D (new_AGEMA_signal_23935), .Q (new_AGEMA_signal_23936) ) ;
    buf_clk new_AGEMA_reg_buffer_11216 ( .C (clk), .D (new_AGEMA_signal_23939), .Q (new_AGEMA_signal_23940) ) ;
    buf_clk new_AGEMA_reg_buffer_11220 ( .C (clk), .D (new_AGEMA_signal_23943), .Q (new_AGEMA_signal_23944) ) ;
    buf_clk new_AGEMA_reg_buffer_11224 ( .C (clk), .D (new_AGEMA_signal_23947), .Q (new_AGEMA_signal_23948) ) ;
    buf_clk new_AGEMA_reg_buffer_11228 ( .C (clk), .D (new_AGEMA_signal_23951), .Q (new_AGEMA_signal_23952) ) ;
    buf_clk new_AGEMA_reg_buffer_11232 ( .C (clk), .D (new_AGEMA_signal_23955), .Q (new_AGEMA_signal_23956) ) ;
    buf_clk new_AGEMA_reg_buffer_11236 ( .C (clk), .D (new_AGEMA_signal_23959), .Q (new_AGEMA_signal_23960) ) ;
    buf_clk new_AGEMA_reg_buffer_11240 ( .C (clk), .D (new_AGEMA_signal_23963), .Q (new_AGEMA_signal_23964) ) ;
    buf_clk new_AGEMA_reg_buffer_11244 ( .C (clk), .D (new_AGEMA_signal_23967), .Q (new_AGEMA_signal_23968) ) ;
    buf_clk new_AGEMA_reg_buffer_11248 ( .C (clk), .D (new_AGEMA_signal_23971), .Q (new_AGEMA_signal_23972) ) ;
    buf_clk new_AGEMA_reg_buffer_11252 ( .C (clk), .D (new_AGEMA_signal_23975), .Q (new_AGEMA_signal_23976) ) ;
    buf_clk new_AGEMA_reg_buffer_11256 ( .C (clk), .D (new_AGEMA_signal_23979), .Q (new_AGEMA_signal_23980) ) ;
    buf_clk new_AGEMA_reg_buffer_11260 ( .C (clk), .D (new_AGEMA_signal_23983), .Q (new_AGEMA_signal_23984) ) ;
    buf_clk new_AGEMA_reg_buffer_11264 ( .C (clk), .D (new_AGEMA_signal_23987), .Q (new_AGEMA_signal_23988) ) ;
    buf_clk new_AGEMA_reg_buffer_11268 ( .C (clk), .D (new_AGEMA_signal_23991), .Q (new_AGEMA_signal_23992) ) ;
    buf_clk new_AGEMA_reg_buffer_11272 ( .C (clk), .D (new_AGEMA_signal_23995), .Q (new_AGEMA_signal_23996) ) ;
    buf_clk new_AGEMA_reg_buffer_11276 ( .C (clk), .D (new_AGEMA_signal_23999), .Q (new_AGEMA_signal_24000) ) ;
    buf_clk new_AGEMA_reg_buffer_11280 ( .C (clk), .D (new_AGEMA_signal_24003), .Q (new_AGEMA_signal_24004) ) ;
    buf_clk new_AGEMA_reg_buffer_11284 ( .C (clk), .D (new_AGEMA_signal_24007), .Q (new_AGEMA_signal_24008) ) ;
    buf_clk new_AGEMA_reg_buffer_11288 ( .C (clk), .D (new_AGEMA_signal_24011), .Q (new_AGEMA_signal_24012) ) ;
    buf_clk new_AGEMA_reg_buffer_11292 ( .C (clk), .D (new_AGEMA_signal_24015), .Q (new_AGEMA_signal_24016) ) ;
    buf_clk new_AGEMA_reg_buffer_11296 ( .C (clk), .D (new_AGEMA_signal_24019), .Q (new_AGEMA_signal_24020) ) ;
    buf_clk new_AGEMA_reg_buffer_11300 ( .C (clk), .D (new_AGEMA_signal_24023), .Q (new_AGEMA_signal_24024) ) ;
    buf_clk new_AGEMA_reg_buffer_11304 ( .C (clk), .D (new_AGEMA_signal_24027), .Q (new_AGEMA_signal_24028) ) ;
    buf_clk new_AGEMA_reg_buffer_11308 ( .C (clk), .D (new_AGEMA_signal_24031), .Q (new_AGEMA_signal_24032) ) ;
    buf_clk new_AGEMA_reg_buffer_11312 ( .C (clk), .D (new_AGEMA_signal_24035), .Q (new_AGEMA_signal_24036) ) ;
    buf_clk new_AGEMA_reg_buffer_11316 ( .C (clk), .D (new_AGEMA_signal_24039), .Q (new_AGEMA_signal_24040) ) ;
    buf_clk new_AGEMA_reg_buffer_11320 ( .C (clk), .D (new_AGEMA_signal_24043), .Q (new_AGEMA_signal_24044) ) ;
    buf_clk new_AGEMA_reg_buffer_11324 ( .C (clk), .D (new_AGEMA_signal_24047), .Q (new_AGEMA_signal_24048) ) ;
    buf_clk new_AGEMA_reg_buffer_11328 ( .C (clk), .D (new_AGEMA_signal_24051), .Q (new_AGEMA_signal_24052) ) ;
    buf_clk new_AGEMA_reg_buffer_11332 ( .C (clk), .D (new_AGEMA_signal_24055), .Q (new_AGEMA_signal_24056) ) ;
    buf_clk new_AGEMA_reg_buffer_11336 ( .C (clk), .D (new_AGEMA_signal_24059), .Q (new_AGEMA_signal_24060) ) ;
    buf_clk new_AGEMA_reg_buffer_11340 ( .C (clk), .D (new_AGEMA_signal_24063), .Q (new_AGEMA_signal_24064) ) ;
    buf_clk new_AGEMA_reg_buffer_11344 ( .C (clk), .D (new_AGEMA_signal_24067), .Q (new_AGEMA_signal_24068) ) ;
    buf_clk new_AGEMA_reg_buffer_11348 ( .C (clk), .D (new_AGEMA_signal_24071), .Q (new_AGEMA_signal_24072) ) ;
    buf_clk new_AGEMA_reg_buffer_11352 ( .C (clk), .D (new_AGEMA_signal_24075), .Q (new_AGEMA_signal_24076) ) ;
    buf_clk new_AGEMA_reg_buffer_11356 ( .C (clk), .D (new_AGEMA_signal_24079), .Q (new_AGEMA_signal_24080) ) ;
    buf_clk new_AGEMA_reg_buffer_11360 ( .C (clk), .D (new_AGEMA_signal_24083), .Q (new_AGEMA_signal_24084) ) ;
    buf_clk new_AGEMA_reg_buffer_11364 ( .C (clk), .D (new_AGEMA_signal_24087), .Q (new_AGEMA_signal_24088) ) ;
    buf_clk new_AGEMA_reg_buffer_11368 ( .C (clk), .D (new_AGEMA_signal_24091), .Q (new_AGEMA_signal_24092) ) ;
    buf_clk new_AGEMA_reg_buffer_11372 ( .C (clk), .D (new_AGEMA_signal_24095), .Q (new_AGEMA_signal_24096) ) ;
    buf_clk new_AGEMA_reg_buffer_11376 ( .C (clk), .D (new_AGEMA_signal_24099), .Q (new_AGEMA_signal_24100) ) ;
    buf_clk new_AGEMA_reg_buffer_11380 ( .C (clk), .D (new_AGEMA_signal_24103), .Q (new_AGEMA_signal_24104) ) ;
    buf_clk new_AGEMA_reg_buffer_11384 ( .C (clk), .D (new_AGEMA_signal_24107), .Q (new_AGEMA_signal_24108) ) ;
    buf_clk new_AGEMA_reg_buffer_11388 ( .C (clk), .D (new_AGEMA_signal_24111), .Q (new_AGEMA_signal_24112) ) ;
    buf_clk new_AGEMA_reg_buffer_11392 ( .C (clk), .D (new_AGEMA_signal_24115), .Q (new_AGEMA_signal_24116) ) ;
    buf_clk new_AGEMA_reg_buffer_11396 ( .C (clk), .D (new_AGEMA_signal_24119), .Q (new_AGEMA_signal_24120) ) ;
    buf_clk new_AGEMA_reg_buffer_11400 ( .C (clk), .D (new_AGEMA_signal_24123), .Q (new_AGEMA_signal_24124) ) ;
    buf_clk new_AGEMA_reg_buffer_11404 ( .C (clk), .D (new_AGEMA_signal_24127), .Q (new_AGEMA_signal_24128) ) ;
    buf_clk new_AGEMA_reg_buffer_11408 ( .C (clk), .D (new_AGEMA_signal_24131), .Q (new_AGEMA_signal_24132) ) ;
    buf_clk new_AGEMA_reg_buffer_11412 ( .C (clk), .D (new_AGEMA_signal_24135), .Q (new_AGEMA_signal_24136) ) ;
    buf_clk new_AGEMA_reg_buffer_11416 ( .C (clk), .D (new_AGEMA_signal_24139), .Q (new_AGEMA_signal_24140) ) ;
    buf_clk new_AGEMA_reg_buffer_11420 ( .C (clk), .D (new_AGEMA_signal_24143), .Q (new_AGEMA_signal_24144) ) ;
    buf_clk new_AGEMA_reg_buffer_11424 ( .C (clk), .D (new_AGEMA_signal_24147), .Q (new_AGEMA_signal_24148) ) ;
    buf_clk new_AGEMA_reg_buffer_11428 ( .C (clk), .D (new_AGEMA_signal_24151), .Q (new_AGEMA_signal_24152) ) ;
    buf_clk new_AGEMA_reg_buffer_11432 ( .C (clk), .D (new_AGEMA_signal_24155), .Q (new_AGEMA_signal_24156) ) ;
    buf_clk new_AGEMA_reg_buffer_11436 ( .C (clk), .D (new_AGEMA_signal_24159), .Q (new_AGEMA_signal_24160) ) ;
    buf_clk new_AGEMA_reg_buffer_11440 ( .C (clk), .D (new_AGEMA_signal_24163), .Q (new_AGEMA_signal_24164) ) ;
    buf_clk new_AGEMA_reg_buffer_11444 ( .C (clk), .D (new_AGEMA_signal_24167), .Q (new_AGEMA_signal_24168) ) ;
    buf_clk new_AGEMA_reg_buffer_11448 ( .C (clk), .D (new_AGEMA_signal_24171), .Q (new_AGEMA_signal_24172) ) ;
    buf_clk new_AGEMA_reg_buffer_11452 ( .C (clk), .D (new_AGEMA_signal_24175), .Q (new_AGEMA_signal_24176) ) ;
    buf_clk new_AGEMA_reg_buffer_11456 ( .C (clk), .D (new_AGEMA_signal_24179), .Q (new_AGEMA_signal_24180) ) ;
    buf_clk new_AGEMA_reg_buffer_11460 ( .C (clk), .D (new_AGEMA_signal_24183), .Q (new_AGEMA_signal_24184) ) ;
    buf_clk new_AGEMA_reg_buffer_11464 ( .C (clk), .D (new_AGEMA_signal_24187), .Q (new_AGEMA_signal_24188) ) ;
    buf_clk new_AGEMA_reg_buffer_11468 ( .C (clk), .D (new_AGEMA_signal_24191), .Q (new_AGEMA_signal_24192) ) ;
    buf_clk new_AGEMA_reg_buffer_11472 ( .C (clk), .D (new_AGEMA_signal_24195), .Q (new_AGEMA_signal_24196) ) ;
    buf_clk new_AGEMA_reg_buffer_11476 ( .C (clk), .D (new_AGEMA_signal_24199), .Q (new_AGEMA_signal_24200) ) ;
    buf_clk new_AGEMA_reg_buffer_11480 ( .C (clk), .D (new_AGEMA_signal_24203), .Q (new_AGEMA_signal_24204) ) ;
    buf_clk new_AGEMA_reg_buffer_11484 ( .C (clk), .D (new_AGEMA_signal_24207), .Q (new_AGEMA_signal_24208) ) ;
    buf_clk new_AGEMA_reg_buffer_11488 ( .C (clk), .D (new_AGEMA_signal_24211), .Q (new_AGEMA_signal_24212) ) ;
    buf_clk new_AGEMA_reg_buffer_11492 ( .C (clk), .D (new_AGEMA_signal_24215), .Q (new_AGEMA_signal_24216) ) ;
    buf_clk new_AGEMA_reg_buffer_11496 ( .C (clk), .D (new_AGEMA_signal_24219), .Q (new_AGEMA_signal_24220) ) ;
    buf_clk new_AGEMA_reg_buffer_11500 ( .C (clk), .D (new_AGEMA_signal_24223), .Q (new_AGEMA_signal_24224) ) ;
    buf_clk new_AGEMA_reg_buffer_11504 ( .C (clk), .D (new_AGEMA_signal_24227), .Q (new_AGEMA_signal_24228) ) ;
    buf_clk new_AGEMA_reg_buffer_11508 ( .C (clk), .D (new_AGEMA_signal_24231), .Q (new_AGEMA_signal_24232) ) ;
    buf_clk new_AGEMA_reg_buffer_11512 ( .C (clk), .D (new_AGEMA_signal_24235), .Q (new_AGEMA_signal_24236) ) ;
    buf_clk new_AGEMA_reg_buffer_11516 ( .C (clk), .D (new_AGEMA_signal_24239), .Q (new_AGEMA_signal_24240) ) ;
    buf_clk new_AGEMA_reg_buffer_11520 ( .C (clk), .D (new_AGEMA_signal_24243), .Q (new_AGEMA_signal_24244) ) ;
    buf_clk new_AGEMA_reg_buffer_11524 ( .C (clk), .D (new_AGEMA_signal_24247), .Q (new_AGEMA_signal_24248) ) ;
    buf_clk new_AGEMA_reg_buffer_11528 ( .C (clk), .D (new_AGEMA_signal_24251), .Q (new_AGEMA_signal_24252) ) ;
    buf_clk new_AGEMA_reg_buffer_11532 ( .C (clk), .D (new_AGEMA_signal_24255), .Q (new_AGEMA_signal_24256) ) ;
    buf_clk new_AGEMA_reg_buffer_11536 ( .C (clk), .D (new_AGEMA_signal_24259), .Q (new_AGEMA_signal_24260) ) ;
    buf_clk new_AGEMA_reg_buffer_11540 ( .C (clk), .D (new_AGEMA_signal_24263), .Q (new_AGEMA_signal_24264) ) ;
    buf_clk new_AGEMA_reg_buffer_11544 ( .C (clk), .D (new_AGEMA_signal_24267), .Q (new_AGEMA_signal_24268) ) ;
    buf_clk new_AGEMA_reg_buffer_11548 ( .C (clk), .D (new_AGEMA_signal_24271), .Q (new_AGEMA_signal_24272) ) ;
    buf_clk new_AGEMA_reg_buffer_11552 ( .C (clk), .D (new_AGEMA_signal_24275), .Q (new_AGEMA_signal_24276) ) ;
    buf_clk new_AGEMA_reg_buffer_11556 ( .C (clk), .D (new_AGEMA_signal_24279), .Q (new_AGEMA_signal_24280) ) ;
    buf_clk new_AGEMA_reg_buffer_11560 ( .C (clk), .D (new_AGEMA_signal_24283), .Q (new_AGEMA_signal_24284) ) ;
    buf_clk new_AGEMA_reg_buffer_11564 ( .C (clk), .D (new_AGEMA_signal_24287), .Q (new_AGEMA_signal_24288) ) ;
    buf_clk new_AGEMA_reg_buffer_11568 ( .C (clk), .D (new_AGEMA_signal_24291), .Q (new_AGEMA_signal_24292) ) ;
    buf_clk new_AGEMA_reg_buffer_11572 ( .C (clk), .D (new_AGEMA_signal_24295), .Q (new_AGEMA_signal_24296) ) ;
    buf_clk new_AGEMA_reg_buffer_11576 ( .C (clk), .D (new_AGEMA_signal_24299), .Q (new_AGEMA_signal_24300) ) ;
    buf_clk new_AGEMA_reg_buffer_11580 ( .C (clk), .D (new_AGEMA_signal_24303), .Q (new_AGEMA_signal_24304) ) ;
    buf_clk new_AGEMA_reg_buffer_11584 ( .C (clk), .D (new_AGEMA_signal_24307), .Q (new_AGEMA_signal_24308) ) ;
    buf_clk new_AGEMA_reg_buffer_11588 ( .C (clk), .D (new_AGEMA_signal_24311), .Q (new_AGEMA_signal_24312) ) ;
    buf_clk new_AGEMA_reg_buffer_11592 ( .C (clk), .D (new_AGEMA_signal_24315), .Q (new_AGEMA_signal_24316) ) ;
    buf_clk new_AGEMA_reg_buffer_11596 ( .C (clk), .D (new_AGEMA_signal_24319), .Q (new_AGEMA_signal_24320) ) ;
    buf_clk new_AGEMA_reg_buffer_11600 ( .C (clk), .D (new_AGEMA_signal_24323), .Q (new_AGEMA_signal_24324) ) ;
    buf_clk new_AGEMA_reg_buffer_11604 ( .C (clk), .D (new_AGEMA_signal_24327), .Q (new_AGEMA_signal_24328) ) ;
    buf_clk new_AGEMA_reg_buffer_11608 ( .C (clk), .D (new_AGEMA_signal_24331), .Q (new_AGEMA_signal_24332) ) ;
    buf_clk new_AGEMA_reg_buffer_11612 ( .C (clk), .D (new_AGEMA_signal_24335), .Q (new_AGEMA_signal_24336) ) ;
    buf_clk new_AGEMA_reg_buffer_11616 ( .C (clk), .D (new_AGEMA_signal_24339), .Q (new_AGEMA_signal_24340) ) ;
    buf_clk new_AGEMA_reg_buffer_11620 ( .C (clk), .D (new_AGEMA_signal_24343), .Q (new_AGEMA_signal_24344) ) ;
    buf_clk new_AGEMA_reg_buffer_11624 ( .C (clk), .D (new_AGEMA_signal_24347), .Q (new_AGEMA_signal_24348) ) ;
    buf_clk new_AGEMA_reg_buffer_11628 ( .C (clk), .D (new_AGEMA_signal_24351), .Q (new_AGEMA_signal_24352) ) ;
    buf_clk new_AGEMA_reg_buffer_11632 ( .C (clk), .D (new_AGEMA_signal_24355), .Q (new_AGEMA_signal_24356) ) ;
    buf_clk new_AGEMA_reg_buffer_11636 ( .C (clk), .D (new_AGEMA_signal_24359), .Q (new_AGEMA_signal_24360) ) ;
    buf_clk new_AGEMA_reg_buffer_11640 ( .C (clk), .D (new_AGEMA_signal_24363), .Q (new_AGEMA_signal_24364) ) ;
    buf_clk new_AGEMA_reg_buffer_11644 ( .C (clk), .D (new_AGEMA_signal_24367), .Q (new_AGEMA_signal_24368) ) ;
    buf_clk new_AGEMA_reg_buffer_11648 ( .C (clk), .D (new_AGEMA_signal_24371), .Q (new_AGEMA_signal_24372) ) ;
    buf_clk new_AGEMA_reg_buffer_11652 ( .C (clk), .D (new_AGEMA_signal_24375), .Q (new_AGEMA_signal_24376) ) ;
    buf_clk new_AGEMA_reg_buffer_11656 ( .C (clk), .D (new_AGEMA_signal_24379), .Q (new_AGEMA_signal_24380) ) ;
    buf_clk new_AGEMA_reg_buffer_11660 ( .C (clk), .D (new_AGEMA_signal_24383), .Q (new_AGEMA_signal_24384) ) ;
    buf_clk new_AGEMA_reg_buffer_11664 ( .C (clk), .D (new_AGEMA_signal_24387), .Q (new_AGEMA_signal_24388) ) ;
    buf_clk new_AGEMA_reg_buffer_11668 ( .C (clk), .D (new_AGEMA_signal_24391), .Q (new_AGEMA_signal_24392) ) ;
    buf_clk new_AGEMA_reg_buffer_11672 ( .C (clk), .D (new_AGEMA_signal_24395), .Q (new_AGEMA_signal_24396) ) ;
    buf_clk new_AGEMA_reg_buffer_11676 ( .C (clk), .D (new_AGEMA_signal_24399), .Q (new_AGEMA_signal_24400) ) ;
    buf_clk new_AGEMA_reg_buffer_11680 ( .C (clk), .D (new_AGEMA_signal_24403), .Q (new_AGEMA_signal_24404) ) ;
    buf_clk new_AGEMA_reg_buffer_11684 ( .C (clk), .D (new_AGEMA_signal_24407), .Q (new_AGEMA_signal_24408) ) ;
    buf_clk new_AGEMA_reg_buffer_11688 ( .C (clk), .D (new_AGEMA_signal_24411), .Q (new_AGEMA_signal_24412) ) ;
    buf_clk new_AGEMA_reg_buffer_11692 ( .C (clk), .D (new_AGEMA_signal_24415), .Q (new_AGEMA_signal_24416) ) ;
    buf_clk new_AGEMA_reg_buffer_11696 ( .C (clk), .D (new_AGEMA_signal_24419), .Q (new_AGEMA_signal_24420) ) ;
    buf_clk new_AGEMA_reg_buffer_11700 ( .C (clk), .D (new_AGEMA_signal_24423), .Q (new_AGEMA_signal_24424) ) ;
    buf_clk new_AGEMA_reg_buffer_11704 ( .C (clk), .D (new_AGEMA_signal_24427), .Q (new_AGEMA_signal_24428) ) ;
    buf_clk new_AGEMA_reg_buffer_11708 ( .C (clk), .D (new_AGEMA_signal_24431), .Q (new_AGEMA_signal_24432) ) ;
    buf_clk new_AGEMA_reg_buffer_11712 ( .C (clk), .D (new_AGEMA_signal_24435), .Q (new_AGEMA_signal_24436) ) ;
    buf_clk new_AGEMA_reg_buffer_11716 ( .C (clk), .D (new_AGEMA_signal_24439), .Q (new_AGEMA_signal_24440) ) ;
    buf_clk new_AGEMA_reg_buffer_11720 ( .C (clk), .D (new_AGEMA_signal_24443), .Q (new_AGEMA_signal_24444) ) ;
    buf_clk new_AGEMA_reg_buffer_11724 ( .C (clk), .D (new_AGEMA_signal_24447), .Q (new_AGEMA_signal_24448) ) ;
    buf_clk new_AGEMA_reg_buffer_11728 ( .C (clk), .D (new_AGEMA_signal_24451), .Q (new_AGEMA_signal_24452) ) ;
    buf_clk new_AGEMA_reg_buffer_11732 ( .C (clk), .D (new_AGEMA_signal_24455), .Q (new_AGEMA_signal_24456) ) ;
    buf_clk new_AGEMA_reg_buffer_11736 ( .C (clk), .D (new_AGEMA_signal_24459), .Q (new_AGEMA_signal_24460) ) ;
    buf_clk new_AGEMA_reg_buffer_11740 ( .C (clk), .D (new_AGEMA_signal_24463), .Q (new_AGEMA_signal_24464) ) ;
    buf_clk new_AGEMA_reg_buffer_11744 ( .C (clk), .D (new_AGEMA_signal_24467), .Q (new_AGEMA_signal_24468) ) ;
    buf_clk new_AGEMA_reg_buffer_11748 ( .C (clk), .D (new_AGEMA_signal_24471), .Q (new_AGEMA_signal_24472) ) ;
    buf_clk new_AGEMA_reg_buffer_11752 ( .C (clk), .D (new_AGEMA_signal_24475), .Q (new_AGEMA_signal_24476) ) ;
    buf_clk new_AGEMA_reg_buffer_11756 ( .C (clk), .D (new_AGEMA_signal_24479), .Q (new_AGEMA_signal_24480) ) ;
    buf_clk new_AGEMA_reg_buffer_11760 ( .C (clk), .D (new_AGEMA_signal_24483), .Q (new_AGEMA_signal_24484) ) ;
    buf_clk new_AGEMA_reg_buffer_11764 ( .C (clk), .D (new_AGEMA_signal_24487), .Q (new_AGEMA_signal_24488) ) ;
    buf_clk new_AGEMA_reg_buffer_11768 ( .C (clk), .D (new_AGEMA_signal_24491), .Q (new_AGEMA_signal_24492) ) ;
    buf_clk new_AGEMA_reg_buffer_11772 ( .C (clk), .D (new_AGEMA_signal_24495), .Q (new_AGEMA_signal_24496) ) ;
    buf_clk new_AGEMA_reg_buffer_11776 ( .C (clk), .D (new_AGEMA_signal_24499), .Q (new_AGEMA_signal_24500) ) ;
    buf_clk new_AGEMA_reg_buffer_11780 ( .C (clk), .D (new_AGEMA_signal_24503), .Q (new_AGEMA_signal_24504) ) ;
    buf_clk new_AGEMA_reg_buffer_11784 ( .C (clk), .D (new_AGEMA_signal_24507), .Q (new_AGEMA_signal_24508) ) ;
    buf_clk new_AGEMA_reg_buffer_11788 ( .C (clk), .D (new_AGEMA_signal_24511), .Q (new_AGEMA_signal_24512) ) ;
    buf_clk new_AGEMA_reg_buffer_11792 ( .C (clk), .D (new_AGEMA_signal_24515), .Q (new_AGEMA_signal_24516) ) ;
    buf_clk new_AGEMA_reg_buffer_11796 ( .C (clk), .D (new_AGEMA_signal_24519), .Q (new_AGEMA_signal_24520) ) ;
    buf_clk new_AGEMA_reg_buffer_11800 ( .C (clk), .D (new_AGEMA_signal_24523), .Q (new_AGEMA_signal_24524) ) ;
    buf_clk new_AGEMA_reg_buffer_11804 ( .C (clk), .D (new_AGEMA_signal_24527), .Q (new_AGEMA_signal_24528) ) ;
    buf_clk new_AGEMA_reg_buffer_11808 ( .C (clk), .D (new_AGEMA_signal_24531), .Q (new_AGEMA_signal_24532) ) ;
    buf_clk new_AGEMA_reg_buffer_11812 ( .C (clk), .D (new_AGEMA_signal_24535), .Q (new_AGEMA_signal_24536) ) ;
    buf_clk new_AGEMA_reg_buffer_11816 ( .C (clk), .D (new_AGEMA_signal_24539), .Q (new_AGEMA_signal_24540) ) ;
    buf_clk new_AGEMA_reg_buffer_11820 ( .C (clk), .D (new_AGEMA_signal_24543), .Q (new_AGEMA_signal_24544) ) ;
    buf_clk new_AGEMA_reg_buffer_11824 ( .C (clk), .D (new_AGEMA_signal_24547), .Q (new_AGEMA_signal_24548) ) ;
    buf_clk new_AGEMA_reg_buffer_11828 ( .C (clk), .D (new_AGEMA_signal_24551), .Q (new_AGEMA_signal_24552) ) ;
    buf_clk new_AGEMA_reg_buffer_11832 ( .C (clk), .D (new_AGEMA_signal_24555), .Q (new_AGEMA_signal_24556) ) ;
    buf_clk new_AGEMA_reg_buffer_11836 ( .C (clk), .D (new_AGEMA_signal_24559), .Q (new_AGEMA_signal_24560) ) ;
    buf_clk new_AGEMA_reg_buffer_11840 ( .C (clk), .D (new_AGEMA_signal_24563), .Q (new_AGEMA_signal_24564) ) ;
    buf_clk new_AGEMA_reg_buffer_11844 ( .C (clk), .D (new_AGEMA_signal_24567), .Q (new_AGEMA_signal_24568) ) ;
    buf_clk new_AGEMA_reg_buffer_11848 ( .C (clk), .D (new_AGEMA_signal_24571), .Q (new_AGEMA_signal_24572) ) ;
    buf_clk new_AGEMA_reg_buffer_11852 ( .C (clk), .D (new_AGEMA_signal_24575), .Q (new_AGEMA_signal_24576) ) ;
    buf_clk new_AGEMA_reg_buffer_11856 ( .C (clk), .D (new_AGEMA_signal_24579), .Q (new_AGEMA_signal_24580) ) ;
    buf_clk new_AGEMA_reg_buffer_11860 ( .C (clk), .D (new_AGEMA_signal_24583), .Q (new_AGEMA_signal_24584) ) ;
    buf_clk new_AGEMA_reg_buffer_11864 ( .C (clk), .D (new_AGEMA_signal_24587), .Q (new_AGEMA_signal_24588) ) ;
    buf_clk new_AGEMA_reg_buffer_11868 ( .C (clk), .D (new_AGEMA_signal_24591), .Q (new_AGEMA_signal_24592) ) ;
    buf_clk new_AGEMA_reg_buffer_11872 ( .C (clk), .D (new_AGEMA_signal_24595), .Q (new_AGEMA_signal_24596) ) ;
    buf_clk new_AGEMA_reg_buffer_11876 ( .C (clk), .D (new_AGEMA_signal_24599), .Q (new_AGEMA_signal_24600) ) ;
    buf_clk new_AGEMA_reg_buffer_11880 ( .C (clk), .D (new_AGEMA_signal_24603), .Q (new_AGEMA_signal_24604) ) ;
    buf_clk new_AGEMA_reg_buffer_11884 ( .C (clk), .D (new_AGEMA_signal_24607), .Q (new_AGEMA_signal_24608) ) ;
    buf_clk new_AGEMA_reg_buffer_11888 ( .C (clk), .D (new_AGEMA_signal_24611), .Q (new_AGEMA_signal_24612) ) ;
    buf_clk new_AGEMA_reg_buffer_11892 ( .C (clk), .D (new_AGEMA_signal_24615), .Q (new_AGEMA_signal_24616) ) ;
    buf_clk new_AGEMA_reg_buffer_11896 ( .C (clk), .D (new_AGEMA_signal_24619), .Q (new_AGEMA_signal_24620) ) ;
    buf_clk new_AGEMA_reg_buffer_11900 ( .C (clk), .D (new_AGEMA_signal_24623), .Q (new_AGEMA_signal_24624) ) ;
    buf_clk new_AGEMA_reg_buffer_11904 ( .C (clk), .D (new_AGEMA_signal_24627), .Q (new_AGEMA_signal_24628) ) ;
    buf_clk new_AGEMA_reg_buffer_11908 ( .C (clk), .D (new_AGEMA_signal_24631), .Q (new_AGEMA_signal_24632) ) ;
    buf_clk new_AGEMA_reg_buffer_11912 ( .C (clk), .D (new_AGEMA_signal_24635), .Q (new_AGEMA_signal_24636) ) ;
    buf_clk new_AGEMA_reg_buffer_11916 ( .C (clk), .D (new_AGEMA_signal_24639), .Q (new_AGEMA_signal_24640) ) ;
    buf_clk new_AGEMA_reg_buffer_11920 ( .C (clk), .D (new_AGEMA_signal_24643), .Q (new_AGEMA_signal_24644) ) ;
    buf_clk new_AGEMA_reg_buffer_11924 ( .C (clk), .D (new_AGEMA_signal_24647), .Q (new_AGEMA_signal_24648) ) ;
    buf_clk new_AGEMA_reg_buffer_11928 ( .C (clk), .D (new_AGEMA_signal_24651), .Q (new_AGEMA_signal_24652) ) ;
    buf_clk new_AGEMA_reg_buffer_11932 ( .C (clk), .D (new_AGEMA_signal_24655), .Q (new_AGEMA_signal_24656) ) ;
    buf_clk new_AGEMA_reg_buffer_11936 ( .C (clk), .D (new_AGEMA_signal_24659), .Q (new_AGEMA_signal_24660) ) ;
    buf_clk new_AGEMA_reg_buffer_11940 ( .C (clk), .D (new_AGEMA_signal_24663), .Q (new_AGEMA_signal_24664) ) ;
    buf_clk new_AGEMA_reg_buffer_11944 ( .C (clk), .D (new_AGEMA_signal_24667), .Q (new_AGEMA_signal_24668) ) ;
    buf_clk new_AGEMA_reg_buffer_11948 ( .C (clk), .D (new_AGEMA_signal_24671), .Q (new_AGEMA_signal_24672) ) ;
    buf_clk new_AGEMA_reg_buffer_11952 ( .C (clk), .D (new_AGEMA_signal_24675), .Q (new_AGEMA_signal_24676) ) ;
    buf_clk new_AGEMA_reg_buffer_11956 ( .C (clk), .D (new_AGEMA_signal_24679), .Q (new_AGEMA_signal_24680) ) ;
    buf_clk new_AGEMA_reg_buffer_11960 ( .C (clk), .D (new_AGEMA_signal_24683), .Q (new_AGEMA_signal_24684) ) ;
    buf_clk new_AGEMA_reg_buffer_11964 ( .C (clk), .D (new_AGEMA_signal_24687), .Q (new_AGEMA_signal_24688) ) ;
    buf_clk new_AGEMA_reg_buffer_11968 ( .C (clk), .D (new_AGEMA_signal_24691), .Q (new_AGEMA_signal_24692) ) ;
    buf_clk new_AGEMA_reg_buffer_11972 ( .C (clk), .D (new_AGEMA_signal_24695), .Q (new_AGEMA_signal_24696) ) ;
    buf_clk new_AGEMA_reg_buffer_11976 ( .C (clk), .D (new_AGEMA_signal_24699), .Q (new_AGEMA_signal_24700) ) ;
    buf_clk new_AGEMA_reg_buffer_11980 ( .C (clk), .D (new_AGEMA_signal_24703), .Q (new_AGEMA_signal_24704) ) ;
    buf_clk new_AGEMA_reg_buffer_11984 ( .C (clk), .D (new_AGEMA_signal_24707), .Q (new_AGEMA_signal_24708) ) ;
    buf_clk new_AGEMA_reg_buffer_11988 ( .C (clk), .D (new_AGEMA_signal_24711), .Q (new_AGEMA_signal_24712) ) ;
    buf_clk new_AGEMA_reg_buffer_11992 ( .C (clk), .D (new_AGEMA_signal_24715), .Q (new_AGEMA_signal_24716) ) ;
    buf_clk new_AGEMA_reg_buffer_11996 ( .C (clk), .D (new_AGEMA_signal_24719), .Q (new_AGEMA_signal_24720) ) ;
    buf_clk new_AGEMA_reg_buffer_12000 ( .C (clk), .D (new_AGEMA_signal_24723), .Q (new_AGEMA_signal_24724) ) ;
    buf_clk new_AGEMA_reg_buffer_12004 ( .C (clk), .D (new_AGEMA_signal_24727), .Q (new_AGEMA_signal_24728) ) ;
    buf_clk new_AGEMA_reg_buffer_12008 ( .C (clk), .D (new_AGEMA_signal_24731), .Q (new_AGEMA_signal_24732) ) ;
    buf_clk new_AGEMA_reg_buffer_12012 ( .C (clk), .D (new_AGEMA_signal_24735), .Q (new_AGEMA_signal_24736) ) ;
    buf_clk new_AGEMA_reg_buffer_12016 ( .C (clk), .D (new_AGEMA_signal_24739), .Q (new_AGEMA_signal_24740) ) ;
    buf_clk new_AGEMA_reg_buffer_12020 ( .C (clk), .D (new_AGEMA_signal_24743), .Q (new_AGEMA_signal_24744) ) ;
    buf_clk new_AGEMA_reg_buffer_12024 ( .C (clk), .D (new_AGEMA_signal_24747), .Q (new_AGEMA_signal_24748) ) ;
    buf_clk new_AGEMA_reg_buffer_12028 ( .C (clk), .D (new_AGEMA_signal_24751), .Q (new_AGEMA_signal_24752) ) ;
    buf_clk new_AGEMA_reg_buffer_12032 ( .C (clk), .D (new_AGEMA_signal_24755), .Q (new_AGEMA_signal_24756) ) ;
    buf_clk new_AGEMA_reg_buffer_12036 ( .C (clk), .D (new_AGEMA_signal_24759), .Q (new_AGEMA_signal_24760) ) ;
    buf_clk new_AGEMA_reg_buffer_12040 ( .C (clk), .D (new_AGEMA_signal_24763), .Q (new_AGEMA_signal_24764) ) ;
    buf_clk new_AGEMA_reg_buffer_12044 ( .C (clk), .D (new_AGEMA_signal_24767), .Q (new_AGEMA_signal_24768) ) ;
    buf_clk new_AGEMA_reg_buffer_12048 ( .C (clk), .D (new_AGEMA_signal_24771), .Q (new_AGEMA_signal_24772) ) ;
    buf_clk new_AGEMA_reg_buffer_12052 ( .C (clk), .D (new_AGEMA_signal_24775), .Q (new_AGEMA_signal_24776) ) ;
    buf_clk new_AGEMA_reg_buffer_12056 ( .C (clk), .D (new_AGEMA_signal_24779), .Q (new_AGEMA_signal_24780) ) ;
    buf_clk new_AGEMA_reg_buffer_12060 ( .C (clk), .D (new_AGEMA_signal_24783), .Q (new_AGEMA_signal_24784) ) ;
    buf_clk new_AGEMA_reg_buffer_12064 ( .C (clk), .D (new_AGEMA_signal_24787), .Q (new_AGEMA_signal_24788) ) ;
    buf_clk new_AGEMA_reg_buffer_12068 ( .C (clk), .D (new_AGEMA_signal_24791), .Q (new_AGEMA_signal_24792) ) ;
    buf_clk new_AGEMA_reg_buffer_12072 ( .C (clk), .D (new_AGEMA_signal_24795), .Q (new_AGEMA_signal_24796) ) ;
    buf_clk new_AGEMA_reg_buffer_12076 ( .C (clk), .D (new_AGEMA_signal_24799), .Q (new_AGEMA_signal_24800) ) ;
    buf_clk new_AGEMA_reg_buffer_12080 ( .C (clk), .D (new_AGEMA_signal_24803), .Q (new_AGEMA_signal_24804) ) ;
    buf_clk new_AGEMA_reg_buffer_12084 ( .C (clk), .D (new_AGEMA_signal_24807), .Q (new_AGEMA_signal_24808) ) ;
    buf_clk new_AGEMA_reg_buffer_12088 ( .C (clk), .D (new_AGEMA_signal_24811), .Q (new_AGEMA_signal_24812) ) ;
    buf_clk new_AGEMA_reg_buffer_12092 ( .C (clk), .D (new_AGEMA_signal_24815), .Q (new_AGEMA_signal_24816) ) ;
    buf_clk new_AGEMA_reg_buffer_12096 ( .C (clk), .D (new_AGEMA_signal_24819), .Q (new_AGEMA_signal_24820) ) ;
    buf_clk new_AGEMA_reg_buffer_12100 ( .C (clk), .D (new_AGEMA_signal_24823), .Q (new_AGEMA_signal_24824) ) ;
    buf_clk new_AGEMA_reg_buffer_12104 ( .C (clk), .D (new_AGEMA_signal_24827), .Q (new_AGEMA_signal_24828) ) ;
    buf_clk new_AGEMA_reg_buffer_12108 ( .C (clk), .D (new_AGEMA_signal_24831), .Q (new_AGEMA_signal_24832) ) ;
    buf_clk new_AGEMA_reg_buffer_12112 ( .C (clk), .D (new_AGEMA_signal_24835), .Q (new_AGEMA_signal_24836) ) ;
    buf_clk new_AGEMA_reg_buffer_12116 ( .C (clk), .D (new_AGEMA_signal_24839), .Q (new_AGEMA_signal_24840) ) ;
    buf_clk new_AGEMA_reg_buffer_12120 ( .C (clk), .D (new_AGEMA_signal_24843), .Q (new_AGEMA_signal_24844) ) ;
    buf_clk new_AGEMA_reg_buffer_12124 ( .C (clk), .D (new_AGEMA_signal_24847), .Q (new_AGEMA_signal_24848) ) ;
    buf_clk new_AGEMA_reg_buffer_12128 ( .C (clk), .D (new_AGEMA_signal_24851), .Q (new_AGEMA_signal_24852) ) ;
    buf_clk new_AGEMA_reg_buffer_12132 ( .C (clk), .D (new_AGEMA_signal_24855), .Q (new_AGEMA_signal_24856) ) ;
    buf_clk new_AGEMA_reg_buffer_12136 ( .C (clk), .D (new_AGEMA_signal_24859), .Q (new_AGEMA_signal_24860) ) ;
    buf_clk new_AGEMA_reg_buffer_12140 ( .C (clk), .D (new_AGEMA_signal_24863), .Q (new_AGEMA_signal_24864) ) ;
    buf_clk new_AGEMA_reg_buffer_12144 ( .C (clk), .D (new_AGEMA_signal_24867), .Q (new_AGEMA_signal_24868) ) ;
    buf_clk new_AGEMA_reg_buffer_12148 ( .C (clk), .D (new_AGEMA_signal_24871), .Q (new_AGEMA_signal_24872) ) ;
    buf_clk new_AGEMA_reg_buffer_12152 ( .C (clk), .D (new_AGEMA_signal_24875), .Q (new_AGEMA_signal_24876) ) ;
    buf_clk new_AGEMA_reg_buffer_12156 ( .C (clk), .D (new_AGEMA_signal_24879), .Q (new_AGEMA_signal_24880) ) ;
    buf_clk new_AGEMA_reg_buffer_12160 ( .C (clk), .D (new_AGEMA_signal_24883), .Q (new_AGEMA_signal_24884) ) ;
    buf_clk new_AGEMA_reg_buffer_12164 ( .C (clk), .D (new_AGEMA_signal_24887), .Q (new_AGEMA_signal_24888) ) ;
    buf_clk new_AGEMA_reg_buffer_12168 ( .C (clk), .D (new_AGEMA_signal_24891), .Q (new_AGEMA_signal_24892) ) ;
    buf_clk new_AGEMA_reg_buffer_12172 ( .C (clk), .D (new_AGEMA_signal_24895), .Q (new_AGEMA_signal_24896) ) ;
    buf_clk new_AGEMA_reg_buffer_12176 ( .C (clk), .D (new_AGEMA_signal_24899), .Q (new_AGEMA_signal_24900) ) ;
    buf_clk new_AGEMA_reg_buffer_12180 ( .C (clk), .D (new_AGEMA_signal_24903), .Q (new_AGEMA_signal_24904) ) ;
    buf_clk new_AGEMA_reg_buffer_12184 ( .C (clk), .D (new_AGEMA_signal_24907), .Q (new_AGEMA_signal_24908) ) ;
    buf_clk new_AGEMA_reg_buffer_12188 ( .C (clk), .D (new_AGEMA_signal_24911), .Q (new_AGEMA_signal_24912) ) ;
    buf_clk new_AGEMA_reg_buffer_12192 ( .C (clk), .D (new_AGEMA_signal_24915), .Q (new_AGEMA_signal_24916) ) ;
    buf_clk new_AGEMA_reg_buffer_12808 ( .C (clk), .D (new_AGEMA_signal_25531), .Q (new_AGEMA_signal_25532) ) ;
    buf_clk new_AGEMA_reg_buffer_12812 ( .C (clk), .D (new_AGEMA_signal_25535), .Q (new_AGEMA_signal_25536) ) ;
    buf_clk new_AGEMA_reg_buffer_12816 ( .C (clk), .D (new_AGEMA_signal_25539), .Q (new_AGEMA_signal_25540) ) ;
    buf_clk new_AGEMA_reg_buffer_12820 ( .C (clk), .D (new_AGEMA_signal_25543), .Q (new_AGEMA_signal_25544) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12320, new_AGEMA_signal_12319, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundInput[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12668, new_AGEMA_signal_12667, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, RoundInput[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundInput[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, RoundInput[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12332, new_AGEMA_signal_12331, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundInput[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5312, new_AGEMA_signal_5311, RoundInput[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundInput[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12680, new_AGEMA_signal_12679, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, RoundInput[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, RoundInput[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12344, new_AGEMA_signal_12343, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundInput[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, RoundInput[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12356, new_AGEMA_signal_12355, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundInput[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, RoundInput[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12692, new_AGEMA_signal_12691, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundInput[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, RoundInput[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundInput[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12368, new_AGEMA_signal_12367, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, RoundInput[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundInput[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12380, new_AGEMA_signal_12379, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, RoundInput[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12704, new_AGEMA_signal_12703, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundInput[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, RoundInput[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12392, new_AGEMA_signal_12391, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, RoundInput[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundInput[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, RoundInput[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12716, new_AGEMA_signal_12715, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundInput[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12404, new_AGEMA_signal_12403, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, RoundInput[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundInput[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12416, new_AGEMA_signal_12415, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundInput[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, RoundInput[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12728, new_AGEMA_signal_12727, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundInput[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, RoundInput[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12428, new_AGEMA_signal_12427, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundInput[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, RoundInput[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundInput[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12440, new_AGEMA_signal_12439, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, RoundInput[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12740, new_AGEMA_signal_12739, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundInput[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, RoundInput[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundInput[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12452, new_AGEMA_signal_12451, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, RoundInput[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundInput[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12752, new_AGEMA_signal_12751, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, RoundInput[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12464, new_AGEMA_signal_12463, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, RoundInput[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundInput[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12476, new_AGEMA_signal_12475, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, RoundInput[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundInput[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12764, new_AGEMA_signal_12763, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, RoundInput[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundInput[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12488, new_AGEMA_signal_12487, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundInput[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, RoundInput[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundInput[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12500, new_AGEMA_signal_12499, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12776, new_AGEMA_signal_12775, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, RoundInput[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundInput[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, RoundInput[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12512, new_AGEMA_signal_12511, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundInput[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, RoundInput[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundInput[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12788, new_AGEMA_signal_12787, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, RoundInput[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundInput[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12524, new_AGEMA_signal_12523, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, RoundInput[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundInput[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12536, new_AGEMA_signal_12535, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, RoundInput[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12800, new_AGEMA_signal_12799, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, RoundInput[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundInput[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12548, new_AGEMA_signal_12547, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, RoundInput[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundInput[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5294, new_AGEMA_signal_5293, RoundInput[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12560, new_AGEMA_signal_12559, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundInput[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12812, new_AGEMA_signal_12811, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, RoundInput[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundInput[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12572, new_AGEMA_signal_12571, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, RoundInput[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundInput[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, RoundInput[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12824, new_AGEMA_signal_12823, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundInput[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12584, new_AGEMA_signal_12583, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, RoundInput[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, RoundInput[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12596, new_AGEMA_signal_12595, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundInput[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, RoundInput[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12836, new_AGEMA_signal_12835, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundInput[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, RoundInput[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12608, new_AGEMA_signal_12607, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundInput[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundInput[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12620, new_AGEMA_signal_12619, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, RoundInput[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12848, new_AGEMA_signal_12847, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundInput[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, RoundInput[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundInput[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12632, new_AGEMA_signal_12631, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[127]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11648, new_AGEMA_signal_11647, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, RoundKey[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, RoundKey[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, RoundKey[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12098, new_AGEMA_signal_12097, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, RoundKey[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, RoundKey[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, RoundKey[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12110, new_AGEMA_signal_12109, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, RoundKey[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, RoundKey[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5248, new_AGEMA_signal_5247, RoundKey[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, RoundKey[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12122, new_AGEMA_signal_12121, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, RoundKey[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, RoundKey[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, RoundKey[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12134, new_AGEMA_signal_12133, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, RoundKey[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, RoundKey[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, RoundKey[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, RoundKey[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12146, new_AGEMA_signal_12145, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, RoundKey[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, RoundKey[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, RoundKey[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12158, new_AGEMA_signal_12157, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, RoundKey[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, RoundKey[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, RoundKey[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12170, new_AGEMA_signal_12169, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, RoundKey[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, RoundKey[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, RoundKey[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, RoundKey[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12644, new_AGEMA_signal_12643, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, RoundKey[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, RoundKey[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, RoundKey[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12656, new_AGEMA_signal_12655, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, RoundKey[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, RoundKey[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, RoundKey[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11660, new_AGEMA_signal_11659, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, RoundKey[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, RoundKey[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, RoundKey[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11672, new_AGEMA_signal_11671, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, RoundKey[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, RoundKey[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, RoundKey[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11684, new_AGEMA_signal_11683, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, RoundKey[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, RoundKey[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, RoundKey[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, RoundKey[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11696, new_AGEMA_signal_11695, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, RoundKey[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, RoundKey[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, RoundKey[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11708, new_AGEMA_signal_11707, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, RoundKey[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, RoundKey[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, RoundKey[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, RoundKey[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11720, new_AGEMA_signal_11719, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, RoundKey[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, RoundKey[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, RoundKey[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11732, new_AGEMA_signal_11731, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, RoundKey[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, RoundKey[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, RoundKey[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11744, new_AGEMA_signal_11743, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, RoundKey[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, RoundKey[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12182, new_AGEMA_signal_12181, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, RoundKey[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, RoundKey[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, RoundKey[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12194, new_AGEMA_signal_12193, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, RoundKey[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, RoundKey[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, RoundKey[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, RoundKey[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, RoundKey[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, RoundKey[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, RoundKey[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, RoundKey[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, RoundKey[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, RoundKey[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, RoundKey[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10784, new_AGEMA_signal_10783, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, RoundKey[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, RoundKey[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, RoundKey[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, RoundKey[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, RoundKey[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, RoundKey[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, RoundKey[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, RoundKey[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, RoundKey[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, RoundKey[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, RoundKey[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5206, new_AGEMA_signal_5205, RoundKey[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5212, new_AGEMA_signal_5211, RoundKey[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5218, new_AGEMA_signal_5217, RoundKey[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11288, new_AGEMA_signal_11287, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5224, new_AGEMA_signal_5223, RoundKey[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, RoundKey[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5236, new_AGEMA_signal_5235, RoundKey[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, RoundKey[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5254, new_AGEMA_signal_5253, RoundKey[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11756, new_AGEMA_signal_11755, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, RoundKey[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, RoundKey[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5272, new_AGEMA_signal_5271, RoundKey[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5278, new_AGEMA_signal_5277, RoundKey[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, RoundKey[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5290, new_AGEMA_signal_5289, RoundKey[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, RoundKey[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10796, new_AGEMA_signal_10795, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5302, new_AGEMA_signal_5301, RoundKey[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5308, new_AGEMA_signal_5307, RoundKey[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, RoundKey[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10808, new_AGEMA_signal_10807, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, RoundKey[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, RoundKey[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, RoundKey[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, RoundKey[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10820, new_AGEMA_signal_10819, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, RoundKey[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, RoundKey[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, RoundKey[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10832, new_AGEMA_signal_10831, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, RoundKey[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, RoundKey[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, RoundKey[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10844, new_AGEMA_signal_10843, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, RoundKey[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, RoundKey[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, RoundKey[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, RoundKey[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10856, new_AGEMA_signal_10855, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, RoundKey[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, RoundKey[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, RoundKey[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10868, new_AGEMA_signal_10867, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, RoundKey[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, RoundKey[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, RoundKey[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11300, new_AGEMA_signal_11299, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, RoundKey[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, RoundKey[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, RoundKey[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11312, new_AGEMA_signal_11311, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, RoundKey[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, RoundKey[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, RoundKey[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_11324, new_AGEMA_signal_11323, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_25532), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_25536), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_25540), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_25544), .Q (RoundCounter[3]), .QN () ) ;
endmodule
