/* modified netlist. Source: module PRESENT in file /PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module PRESENT_HPC2_BDDcudd_ClockGating_d1 (data_in_s0, key_s0, clk, reset, data_in_s1, key_s1, Fresh, data_out_s0, done, data_out_s1, Synch);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [21:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    output Synch ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_443 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_885 ;
    wire signal_888 ;
    wire signal_891 ;
    wire signal_894 ;
    wire signal_897 ;
    wire signal_900 ;
    wire signal_903 ;
    wire signal_906 ;
    wire signal_909 ;
    wire signal_912 ;
    wire signal_915 ;
    wire signal_918 ;
    wire signal_921 ;
    wire signal_924 ;
    wire signal_927 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_935 ;
    wire signal_938 ;
    wire signal_941 ;
    wire signal_944 ;
    wire signal_947 ;
    wire signal_950 ;
    wire signal_953 ;
    wire signal_956 ;
    wire signal_959 ;
    wire signal_962 ;
    wire signal_965 ;
    wire signal_968 ;
    wire signal_971 ;
    wire signal_974 ;
    wire signal_977 ;
    wire signal_979 ;
    wire signal_982 ;
    wire signal_985 ;
    wire signal_988 ;
    wire signal_991 ;
    wire signal_994 ;
    wire signal_997 ;
    wire signal_1000 ;
    wire signal_1003 ;
    wire signal_1006 ;
    wire signal_1009 ;
    wire signal_1012 ;
    wire signal_1015 ;
    wire signal_1018 ;
    wire signal_1021 ;
    wire signal_1024 ;
    wire signal_1026 ;
    wire signal_1029 ;
    wire signal_1032 ;
    wire signal_1035 ;
    wire signal_1038 ;
    wire signal_1041 ;
    wire signal_1044 ;
    wire signal_1047 ;
    wire signal_1050 ;
    wire signal_1053 ;
    wire signal_1056 ;
    wire signal_1059 ;
    wire signal_1062 ;
    wire signal_1065 ;
    wire signal_1068 ;
    wire signal_1071 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1297 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1470 ;
    wire signal_1472 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1512 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_0 ( .a ({signal_874, signal_474}), .b ({data_out_s1[60], data_out_s0[60]}), .c ({signal_876, signal_485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_1 ( .a ({signal_877, signal_473}), .b ({data_out_s1[61], data_out_s0[61]}), .c ({signal_879, signal_484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_2 ( .a ({signal_880, signal_472}), .b ({data_out_s1[62], data_out_s0[62]}), .c ({signal_882, signal_483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3 ( .a ({signal_883, signal_471}), .b ({data_out_s1[63], data_out_s0[63]}), .c ({signal_885, signal_482}) ) ;
    NOR2_X1 cell_4 ( .A1 (reset), .A2 (signal_220), .ZN (signal_236) ) ;
    NOR2_X1 cell_5 ( .A1 (signal_221), .A2 (done), .ZN (signal_220) ) ;
    NOR2_X1 cell_6 ( .A1 (reset), .A2 (signal_222), .ZN (signal_233) ) ;
    NOR2_X1 cell_7 ( .A1 (signal_235), .A2 (signal_223), .ZN (signal_222) ) ;
    NOR2_X1 cell_8 ( .A1 (signal_224), .A2 (signal_225), .ZN (signal_223) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_459), .A2 (signal_461), .ZN (signal_225) ) ;
    OR2_X1 cell_10 ( .A1 (signal_226), .A2 (signal_227), .ZN (signal_224) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_462), .A2 (signal_458), .ZN (signal_227) ) ;
    NAND2_X1 cell_12 ( .A1 (signal_460), .A2 (signal_234), .ZN (signal_226) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_237), .A2 (signal_232), .ZN (done) ) ;
    AND2_X1 cell_14 ( .A1 (signal_221), .A2 (signal_232), .ZN (signal_239) ) ;
    AND2_X1 cell_15 ( .A1 (signal_487), .A2 (signal_228), .ZN (signal_221) ) ;
    NOR2_X1 cell_16 ( .A1 (signal_229), .A2 (signal_230), .ZN (signal_228) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_488), .A2 (signal_489), .ZN (signal_230) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_237), .A2 (signal_486), .ZN (signal_229) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_234), .A2 (signal_232), .ZN (signal_219) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_235), .A2 (signal_237), .ZN (signal_217) ) ;
    NOR2_X1 cell_21 ( .A1 (reset), .A2 (signal_217), .ZN (signal_238) ) ;
    INV_X1 cell_22 ( .A (reset), .ZN (signal_231) ) ;
    INV_X1 cell_23 ( .A (signal_238), .ZN (signal_218) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_240), .A2 (signal_241), .ZN (signal_266) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_242), .A2 (signal_461), .ZN (signal_241) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_243), .A2 (signal_265), .ZN (signal_240) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_244), .A2 (signal_462), .ZN (signal_243) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_245), .A2 (signal_246), .ZN (signal_269) ) ;
    NAND2_X1 cell_29 ( .A1 (signal_247), .A2 (signal_462), .ZN (signal_246) ) ;
    MUX2_X1 cell_30 ( .S (signal_263), .A (signal_248), .B (signal_249), .Z (signal_270) ) ;
    NAND2_X1 cell_31 ( .A1 (signal_242), .A2 (signal_250), .ZN (signal_248) ) ;
    NAND2_X1 cell_32 ( .A1 (signal_244), .A2 (signal_265), .ZN (signal_250) ) ;
    NOR2_X1 cell_33 ( .A1 (signal_251), .A2 (signal_247), .ZN (signal_242) ) ;
    NOR2_X1 cell_34 ( .A1 (signal_239), .A2 (signal_262), .ZN (signal_247) ) ;
    INV_X1 cell_35 ( .A (signal_245), .ZN (signal_251) ) ;
    NAND2_X1 cell_36 ( .A1 (signal_244), .A2 (signal_264), .ZN (signal_245) ) ;
    MUX2_X1 cell_37 ( .S (signal_458), .A (signal_252), .B (signal_253), .Z (signal_271) ) ;
    NAND2_X1 cell_38 ( .A1 (signal_254), .A2 (signal_255), .ZN (signal_253) ) ;
    NAND2_X1 cell_39 ( .A1 (signal_244), .A2 (signal_267), .ZN (signal_254) ) ;
    INV_X1 cell_40 ( .A (signal_256), .ZN (signal_244) ) ;
    NOR2_X1 cell_41 ( .A1 (signal_267), .A2 (signal_257), .ZN (signal_252) ) ;
    INV_X1 cell_42 ( .A (signal_258), .ZN (signal_268) ) ;
    MUX2_X1 cell_43 ( .S (signal_267), .A (signal_255), .B (signal_257), .Z (signal_258) ) ;
    NAND2_X1 cell_44 ( .A1 (signal_460), .A2 (signal_249), .ZN (signal_257) ) ;
    NOR2_X1 cell_45 ( .A1 (signal_256), .A2 (signal_259), .ZN (signal_249) ) ;
    NAND2_X1 cell_46 ( .A1 (signal_239), .A2 (signal_231), .ZN (signal_256) ) ;
    NAND2_X1 cell_47 ( .A1 (signal_231), .A2 (signal_260), .ZN (signal_255) ) ;
    NAND2_X1 cell_48 ( .A1 (signal_239), .A2 (signal_261), .ZN (signal_260) ) ;
    NOR2_X1 cell_49 ( .A1 (signal_263), .A2 (signal_259), .ZN (signal_261) ) ;
    OR2_X1 cell_50 ( .A1 (signal_265), .A2 (signal_264), .ZN (signal_259) ) ;
    INV_X1 cell_51 ( .A (signal_231), .ZN (signal_262) ) ;
    INV_X1 cell_54 ( .A (signal_460), .ZN (signal_263) ) ;
    INV_X1 cell_56 ( .A (signal_462), .ZN (signal_264) ) ;
    INV_X1 cell_58 ( .A (signal_459), .ZN (signal_267) ) ;
    INV_X1 cell_60 ( .A (signal_265), .ZN (signal_461) ) ;
    NOR2_X1 cell_62 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_284) ) ;
    XNOR2_X1 cell_63 ( .A (signal_237), .B (signal_489), .ZN (signal_273) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_274), .A2 (signal_275), .ZN (signal_282) ) ;
    XOR2_X1 cell_65 ( .A (signal_488), .B (signal_276), .Z (signal_275) ) ;
    NOR2_X1 cell_66 ( .A1 (signal_274), .A2 (signal_277), .ZN (signal_283) ) ;
    XOR2_X1 cell_67 ( .A (signal_486), .B (signal_278), .Z (signal_277) ) ;
    NAND2_X1 cell_68 ( .A1 (signal_279), .A2 (signal_487), .ZN (signal_278) ) ;
    NOR2_X1 cell_69 ( .A1 (signal_280), .A2 (signal_274), .ZN (signal_285) ) ;
    INV_X1 cell_70 ( .A (signal_238), .ZN (signal_274) ) ;
    XNOR2_X1 cell_71 ( .A (signal_279), .B (signal_487), .ZN (signal_280) ) ;
    NOR2_X1 cell_72 ( .A1 (signal_281), .A2 (signal_276), .ZN (signal_279) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_237), .A2 (signal_489), .ZN (signal_276) ) ;
    INV_X1 cell_80 ( .A (signal_488), .ZN (signal_281) ) ;
    INV_X1 cell_82 ( .A (signal_234), .ZN (signal_237) ) ;
    INV_X1 cell_84 ( .A (signal_235), .ZN (signal_232) ) ;
    INV_X1 cell_86 ( .A (signal_289), .ZN (signal_290) ) ;
    INV_X1 cell_87 ( .A (signal_289), .ZN (signal_291) ) ;
    INV_X1 cell_88 ( .A (signal_218), .ZN (signal_289) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_109 ( .s (signal_218), .b ({data_out_s1[0], data_out_s0[0]}), .a ({signal_900, signal_549}), .c ({signal_1315, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_110 ( .s (signal_218), .b ({data_out_s1[1], data_out_s0[1]}), .a ({signal_903, signal_548}), .c ({signal_1316, signal_560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_111 ( .s (signal_218), .b ({data_out_s1[2], data_out_s0[2]}), .a ({signal_906, signal_547}), .c ({signal_1317, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_112 ( .s (signal_218), .b ({data_out_s1[3], data_out_s0[3]}), .a ({signal_909, signal_546}), .c ({signal_1318, signal_558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_121 ( .s (signal_290), .b ({data_out_s1[4], data_out_s0[4]}), .a ({signal_912, signal_545}), .c ({signal_1341, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_122 ( .s (signal_290), .b ({data_out_s1[5], data_out_s0[5]}), .a ({signal_915, signal_544}), .c ({signal_1342, signal_564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_123 ( .s (signal_290), .b ({data_out_s1[6], data_out_s0[6]}), .a ({signal_918, signal_543}), .c ({signal_1343, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_124 ( .s (signal_290), .b ({data_out_s1[7], data_out_s0[7]}), .a ({signal_921, signal_542}), .c ({signal_1344, signal_562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_133 ( .s (signal_290), .b ({data_out_s1[8], data_out_s0[8]}), .a ({signal_924, signal_541}), .c ({signal_1345, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_134 ( .s (signal_290), .b ({data_out_s1[9], data_out_s0[9]}), .a ({signal_927, signal_540}), .c ({signal_1346, signal_568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_135 ( .s (signal_290), .b ({data_out_s1[10], data_out_s0[10]}), .a ({signal_930, signal_539}), .c ({signal_1347, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_136 ( .s (signal_290), .b ({data_out_s1[11], data_out_s0[11]}), .a ({signal_932, signal_538}), .c ({signal_1348, signal_566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_145 ( .s (signal_290), .b ({data_out_s1[12], data_out_s0[12]}), .a ({signal_935, signal_537}), .c ({signal_1349, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_146 ( .s (signal_290), .b ({data_out_s1[13], data_out_s0[13]}), .a ({signal_938, signal_536}), .c ({signal_1350, signal_572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_147 ( .s (signal_290), .b ({data_out_s1[14], data_out_s0[14]}), .a ({signal_941, signal_535}), .c ({signal_1351, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_148 ( .s (signal_290), .b ({data_out_s1[15], data_out_s0[15]}), .a ({signal_944, signal_534}), .c ({signal_1352, signal_570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_157 ( .s (signal_290), .b ({data_out_s1[16], data_out_s0[16]}), .a ({signal_947, signal_533}), .c ({signal_1353, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_158 ( .s (signal_290), .b ({data_out_s1[17], data_out_s0[17]}), .a ({signal_950, signal_532}), .c ({signal_1354, signal_576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_159 ( .s (signal_290), .b ({data_out_s1[18], data_out_s0[18]}), .a ({signal_953, signal_531}), .c ({signal_1355, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_160 ( .s (signal_290), .b ({data_out_s1[19], data_out_s0[19]}), .a ({signal_956, signal_530}), .c ({signal_1356, signal_574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_169 ( .s (signal_290), .b ({data_out_s1[20], data_out_s0[20]}), .a ({signal_959, signal_529}), .c ({signal_1357, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_170 ( .s (signal_290), .b ({data_out_s1[21], data_out_s0[21]}), .a ({signal_962, signal_528}), .c ({signal_1358, signal_580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_171 ( .s (signal_290), .b ({data_out_s1[22], data_out_s0[22]}), .a ({signal_965, signal_527}), .c ({signal_1359, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_172 ( .s (signal_290), .b ({data_out_s1[23], data_out_s0[23]}), .a ({signal_968, signal_526}), .c ({signal_1360, signal_578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_181 ( .s (signal_290), .b ({data_out_s1[24], data_out_s0[24]}), .a ({signal_971, signal_525}), .c ({signal_1361, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_182 ( .s (signal_290), .b ({data_out_s1[25], data_out_s0[25]}), .a ({signal_974, signal_524}), .c ({signal_1362, signal_584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_183 ( .s (signal_290), .b ({data_out_s1[26], data_out_s0[26]}), .a ({signal_977, signal_523}), .c ({signal_1363, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_184 ( .s (signal_290), .b ({data_out_s1[27], data_out_s0[27]}), .a ({signal_979, signal_522}), .c ({signal_1364, signal_582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_193 ( .s (signal_290), .b ({data_out_s1[28], data_out_s0[28]}), .a ({signal_982, signal_521}), .c ({signal_1365, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_194 ( .s (signal_290), .b ({data_out_s1[29], data_out_s0[29]}), .a ({signal_985, signal_520}), .c ({signal_1366, signal_588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_195 ( .s (signal_290), .b ({data_out_s1[30], data_out_s0[30]}), .a ({signal_988, signal_519}), .c ({signal_1367, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_196 ( .s (signal_290), .b ({data_out_s1[31], data_out_s0[31]}), .a ({signal_991, signal_518}), .c ({signal_1368, signal_586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_205 ( .s (signal_291), .b ({data_out_s1[32], data_out_s0[32]}), .a ({signal_994, signal_517}), .c ({signal_1369, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_206 ( .s (signal_291), .b ({data_out_s1[33], data_out_s0[33]}), .a ({signal_997, signal_516}), .c ({signal_1370, signal_592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_207 ( .s (signal_291), .b ({data_out_s1[34], data_out_s0[34]}), .a ({signal_1000, signal_515}), .c ({signal_1371, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_208 ( .s (signal_291), .b ({data_out_s1[35], data_out_s0[35]}), .a ({signal_1003, signal_514}), .c ({signal_1372, signal_590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_217 ( .s (signal_291), .b ({data_out_s1[36], data_out_s0[36]}), .a ({signal_1006, signal_513}), .c ({signal_1373, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_218 ( .s (signal_291), .b ({data_out_s1[37], data_out_s0[37]}), .a ({signal_1009, signal_512}), .c ({signal_1374, signal_596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_219 ( .s (signal_291), .b ({data_out_s1[38], data_out_s0[38]}), .a ({signal_1012, signal_511}), .c ({signal_1375, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_220 ( .s (signal_291), .b ({data_out_s1[39], data_out_s0[39]}), .a ({signal_1015, signal_510}), .c ({signal_1376, signal_594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_229 ( .s (signal_291), .b ({data_out_s1[40], data_out_s0[40]}), .a ({signal_1018, signal_509}), .c ({signal_1377, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_230 ( .s (signal_291), .b ({data_out_s1[41], data_out_s0[41]}), .a ({signal_1021, signal_508}), .c ({signal_1378, signal_600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_231 ( .s (signal_291), .b ({data_out_s1[42], data_out_s0[42]}), .a ({signal_1024, signal_507}), .c ({signal_1379, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_232 ( .s (signal_291), .b ({data_out_s1[43], data_out_s0[43]}), .a ({signal_1026, signal_506}), .c ({signal_1380, signal_598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_241 ( .s (signal_291), .b ({data_out_s1[44], data_out_s0[44]}), .a ({signal_1029, signal_505}), .c ({signal_1381, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_242 ( .s (signal_291), .b ({data_out_s1[45], data_out_s0[45]}), .a ({signal_1032, signal_504}), .c ({signal_1382, signal_604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_243 ( .s (signal_291), .b ({data_out_s1[46], data_out_s0[46]}), .a ({signal_1035, signal_503}), .c ({signal_1383, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_244 ( .s (signal_291), .b ({data_out_s1[47], data_out_s0[47]}), .a ({signal_1038, signal_502}), .c ({signal_1384, signal_602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_253 ( .s (signal_291), .b ({data_out_s1[48], data_out_s0[48]}), .a ({signal_1041, signal_501}), .c ({signal_1385, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_254 ( .s (signal_291), .b ({data_out_s1[49], data_out_s0[49]}), .a ({signal_1044, signal_500}), .c ({signal_1386, signal_608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_255 ( .s (signal_291), .b ({data_out_s1[50], data_out_s0[50]}), .a ({signal_1047, signal_499}), .c ({signal_1387, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_256 ( .s (signal_291), .b ({data_out_s1[51], data_out_s0[51]}), .a ({signal_1050, signal_498}), .c ({signal_1388, signal_606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_265 ( .s (signal_291), .b ({data_out_s1[52], data_out_s0[52]}), .a ({signal_1053, signal_497}), .c ({signal_1389, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_266 ( .s (signal_291), .b ({data_out_s1[53], data_out_s0[53]}), .a ({signal_1056, signal_496}), .c ({signal_1390, signal_612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_267 ( .s (signal_291), .b ({data_out_s1[54], data_out_s0[54]}), .a ({signal_1059, signal_495}), .c ({signal_1391, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_268 ( .s (signal_291), .b ({data_out_s1[55], data_out_s0[55]}), .a ({signal_1062, signal_494}), .c ({signal_1392, signal_610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_277 ( .s (signal_291), .b ({data_out_s1[56], data_out_s0[56]}), .a ({signal_1065, signal_493}), .c ({signal_1393, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_278 ( .s (signal_291), .b ({data_out_s1[57], data_out_s0[57]}), .a ({signal_1068, signal_492}), .c ({signal_1394, signal_616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_279 ( .s (signal_291), .b ({data_out_s1[58], data_out_s0[58]}), .a ({signal_1071, signal_491}), .c ({signal_1395, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_280 ( .s (signal_291), .b ({data_out_s1[59], data_out_s0[59]}), .a ({signal_1073, signal_490}), .c ({signal_1396, signal_614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_281 ( .s (reset), .b ({data_out_s1[0], data_out_s0[0]}), .a ({data_in_s1[0], data_in_s0[0]}), .c ({signal_888, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_282 ( .s (reset), .b ({data_out_s1[4], data_out_s0[4]}), .a ({data_in_s1[1], data_in_s0[1]}), .c ({signal_891, signal_552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_283 ( .s (reset), .b ({data_out_s1[8], data_out_s0[8]}), .a ({data_in_s1[2], data_in_s0[2]}), .c ({signal_894, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_284 ( .s (reset), .b ({data_out_s1[12], data_out_s0[12]}), .a ({data_in_s1[3], data_in_s0[3]}), .c ({signal_897, signal_550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_285 ( .s (reset), .b ({data_out_s1[16], data_out_s0[16]}), .a ({data_in_s1[4], data_in_s0[4]}), .c ({signal_900, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_286 ( .s (reset), .b ({data_out_s1[20], data_out_s0[20]}), .a ({data_in_s1[5], data_in_s0[5]}), .c ({signal_903, signal_548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_287 ( .s (reset), .b ({data_out_s1[24], data_out_s0[24]}), .a ({data_in_s1[6], data_in_s0[6]}), .c ({signal_906, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_288 ( .s (reset), .b ({data_out_s1[28], data_out_s0[28]}), .a ({data_in_s1[7], data_in_s0[7]}), .c ({signal_909, signal_546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_289 ( .s (reset), .b ({data_out_s1[32], data_out_s0[32]}), .a ({data_in_s1[8], data_in_s0[8]}), .c ({signal_912, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_290 ( .s (reset), .b ({data_out_s1[36], data_out_s0[36]}), .a ({data_in_s1[9], data_in_s0[9]}), .c ({signal_915, signal_544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_291 ( .s (reset), .b ({data_out_s1[40], data_out_s0[40]}), .a ({data_in_s1[10], data_in_s0[10]}), .c ({signal_918, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_292 ( .s (reset), .b ({data_out_s1[44], data_out_s0[44]}), .a ({data_in_s1[11], data_in_s0[11]}), .c ({signal_921, signal_542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_293 ( .s (reset), .b ({data_out_s1[48], data_out_s0[48]}), .a ({data_in_s1[12], data_in_s0[12]}), .c ({signal_924, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_294 ( .s (reset), .b ({data_out_s1[52], data_out_s0[52]}), .a ({data_in_s1[13], data_in_s0[13]}), .c ({signal_927, signal_540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_295 ( .s (reset), .b ({data_out_s1[56], data_out_s0[56]}), .a ({data_in_s1[14], data_in_s0[14]}), .c ({signal_930, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_296 ( .s (reset), .b ({data_out_s1[60], data_out_s0[60]}), .a ({data_in_s1[15], data_in_s0[15]}), .c ({signal_932, signal_538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_297 ( .s (reset), .b ({data_out_s1[1], data_out_s0[1]}), .a ({data_in_s1[16], data_in_s0[16]}), .c ({signal_935, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_298 ( .s (reset), .b ({data_out_s1[5], data_out_s0[5]}), .a ({data_in_s1[17], data_in_s0[17]}), .c ({signal_938, signal_536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_299 ( .s (reset), .b ({data_out_s1[9], data_out_s0[9]}), .a ({data_in_s1[18], data_in_s0[18]}), .c ({signal_941, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_300 ( .s (reset), .b ({data_out_s1[13], data_out_s0[13]}), .a ({data_in_s1[19], data_in_s0[19]}), .c ({signal_944, signal_534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_301 ( .s (reset), .b ({data_out_s1[17], data_out_s0[17]}), .a ({data_in_s1[20], data_in_s0[20]}), .c ({signal_947, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_302 ( .s (reset), .b ({data_out_s1[21], data_out_s0[21]}), .a ({data_in_s1[21], data_in_s0[21]}), .c ({signal_950, signal_532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_303 ( .s (reset), .b ({data_out_s1[25], data_out_s0[25]}), .a ({data_in_s1[22], data_in_s0[22]}), .c ({signal_953, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_304 ( .s (reset), .b ({data_out_s1[29], data_out_s0[29]}), .a ({data_in_s1[23], data_in_s0[23]}), .c ({signal_956, signal_530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_305 ( .s (reset), .b ({data_out_s1[33], data_out_s0[33]}), .a ({data_in_s1[24], data_in_s0[24]}), .c ({signal_959, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_306 ( .s (reset), .b ({data_out_s1[37], data_out_s0[37]}), .a ({data_in_s1[25], data_in_s0[25]}), .c ({signal_962, signal_528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_307 ( .s (reset), .b ({data_out_s1[41], data_out_s0[41]}), .a ({data_in_s1[26], data_in_s0[26]}), .c ({signal_965, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_308 ( .s (reset), .b ({data_out_s1[45], data_out_s0[45]}), .a ({data_in_s1[27], data_in_s0[27]}), .c ({signal_968, signal_526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_309 ( .s (reset), .b ({data_out_s1[49], data_out_s0[49]}), .a ({data_in_s1[28], data_in_s0[28]}), .c ({signal_971, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_310 ( .s (reset), .b ({data_out_s1[53], data_out_s0[53]}), .a ({data_in_s1[29], data_in_s0[29]}), .c ({signal_974, signal_524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_311 ( .s (reset), .b ({data_out_s1[57], data_out_s0[57]}), .a ({data_in_s1[30], data_in_s0[30]}), .c ({signal_977, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_312 ( .s (reset), .b ({data_out_s1[61], data_out_s0[61]}), .a ({data_in_s1[31], data_in_s0[31]}), .c ({signal_979, signal_522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_313 ( .s (reset), .b ({data_out_s1[2], data_out_s0[2]}), .a ({data_in_s1[32], data_in_s0[32]}), .c ({signal_982, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_314 ( .s (reset), .b ({data_out_s1[6], data_out_s0[6]}), .a ({data_in_s1[33], data_in_s0[33]}), .c ({signal_985, signal_520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_315 ( .s (reset), .b ({data_out_s1[10], data_out_s0[10]}), .a ({data_in_s1[34], data_in_s0[34]}), .c ({signal_988, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_316 ( .s (reset), .b ({data_out_s1[14], data_out_s0[14]}), .a ({data_in_s1[35], data_in_s0[35]}), .c ({signal_991, signal_518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_317 ( .s (reset), .b ({data_out_s1[18], data_out_s0[18]}), .a ({data_in_s1[36], data_in_s0[36]}), .c ({signal_994, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_318 ( .s (reset), .b ({data_out_s1[22], data_out_s0[22]}), .a ({data_in_s1[37], data_in_s0[37]}), .c ({signal_997, signal_516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_319 ( .s (reset), .b ({data_out_s1[26], data_out_s0[26]}), .a ({data_in_s1[38], data_in_s0[38]}), .c ({signal_1000, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_320 ( .s (reset), .b ({data_out_s1[30], data_out_s0[30]}), .a ({data_in_s1[39], data_in_s0[39]}), .c ({signal_1003, signal_514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_321 ( .s (reset), .b ({data_out_s1[34], data_out_s0[34]}), .a ({data_in_s1[40], data_in_s0[40]}), .c ({signal_1006, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_322 ( .s (reset), .b ({data_out_s1[38], data_out_s0[38]}), .a ({data_in_s1[41], data_in_s0[41]}), .c ({signal_1009, signal_512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_323 ( .s (reset), .b ({data_out_s1[42], data_out_s0[42]}), .a ({data_in_s1[42], data_in_s0[42]}), .c ({signal_1012, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_324 ( .s (reset), .b ({data_out_s1[46], data_out_s0[46]}), .a ({data_in_s1[43], data_in_s0[43]}), .c ({signal_1015, signal_510}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_325 ( .s (reset), .b ({data_out_s1[50], data_out_s0[50]}), .a ({data_in_s1[44], data_in_s0[44]}), .c ({signal_1018, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_326 ( .s (reset), .b ({data_out_s1[54], data_out_s0[54]}), .a ({data_in_s1[45], data_in_s0[45]}), .c ({signal_1021, signal_508}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_327 ( .s (reset), .b ({data_out_s1[58], data_out_s0[58]}), .a ({data_in_s1[46], data_in_s0[46]}), .c ({signal_1024, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_328 ( .s (reset), .b ({data_out_s1[62], data_out_s0[62]}), .a ({data_in_s1[47], data_in_s0[47]}), .c ({signal_1026, signal_506}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_329 ( .s (reset), .b ({data_out_s1[3], data_out_s0[3]}), .a ({data_in_s1[48], data_in_s0[48]}), .c ({signal_1029, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_330 ( .s (reset), .b ({data_out_s1[7], data_out_s0[7]}), .a ({data_in_s1[49], data_in_s0[49]}), .c ({signal_1032, signal_504}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_331 ( .s (reset), .b ({data_out_s1[11], data_out_s0[11]}), .a ({data_in_s1[50], data_in_s0[50]}), .c ({signal_1035, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_332 ( .s (reset), .b ({data_out_s1[15], data_out_s0[15]}), .a ({data_in_s1[51], data_in_s0[51]}), .c ({signal_1038, signal_502}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_333 ( .s (reset), .b ({data_out_s1[19], data_out_s0[19]}), .a ({data_in_s1[52], data_in_s0[52]}), .c ({signal_1041, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_334 ( .s (reset), .b ({data_out_s1[23], data_out_s0[23]}), .a ({data_in_s1[53], data_in_s0[53]}), .c ({signal_1044, signal_500}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_335 ( .s (reset), .b ({data_out_s1[27], data_out_s0[27]}), .a ({data_in_s1[54], data_in_s0[54]}), .c ({signal_1047, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_336 ( .s (reset), .b ({data_out_s1[31], data_out_s0[31]}), .a ({data_in_s1[55], data_in_s0[55]}), .c ({signal_1050, signal_498}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_337 ( .s (reset), .b ({data_out_s1[35], data_out_s0[35]}), .a ({data_in_s1[56], data_in_s0[56]}), .c ({signal_1053, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_338 ( .s (reset), .b ({data_out_s1[39], data_out_s0[39]}), .a ({data_in_s1[57], data_in_s0[57]}), .c ({signal_1056, signal_496}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_339 ( .s (reset), .b ({data_out_s1[43], data_out_s0[43]}), .a ({data_in_s1[58], data_in_s0[58]}), .c ({signal_1059, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_340 ( .s (reset), .b ({data_out_s1[47], data_out_s0[47]}), .a ({data_in_s1[59], data_in_s0[59]}), .c ({signal_1062, signal_494}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_341 ( .s (reset), .b ({data_out_s1[51], data_out_s0[51]}), .a ({data_in_s1[60], data_in_s0[60]}), .c ({signal_1065, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_342 ( .s (reset), .b ({data_out_s1[55], data_out_s0[55]}), .a ({data_in_s1[61], data_in_s0[61]}), .c ({signal_1068, signal_492}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_343 ( .s (reset), .b ({data_out_s1[59], data_out_s0[59]}), .a ({data_in_s1[62], data_in_s0[62]}), .c ({signal_1071, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_344 ( .s (reset), .b ({data_out_s1[63], data_out_s0[63]}), .a ({data_in_s1[63], data_in_s0[63]}), .c ({signal_1073, signal_490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_345 ( .a ({1'b0, signal_458}), .b ({signal_1074, signal_676}), .c ({signal_1075, signal_618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_346 ( .a ({1'b0, signal_459}), .b ({signal_1076, signal_677}), .c ({signal_1077, signal_619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_347 ( .a ({1'b0, signal_460}), .b ({signal_1078, signal_678}), .c ({signal_1079, signal_620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_348 ( .a ({1'b0, signal_461}), .b ({signal_1292, signal_679}), .c ({signal_1293, signal_621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_349 ( .a ({1'b0, signal_462}), .b ({signal_1080, signal_680}), .c ({signal_1081, signal_622}) ) ;
    INV_X1 cell_350 ( .A (signal_356), .ZN (signal_358) ) ;
    INV_X1 cell_351 ( .A (signal_356), .ZN (signal_357) ) ;
    INV_X1 cell_352 ( .A (signal_218), .ZN (signal_356) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_361 ( .s (signal_357), .b ({signal_874, signal_474}), .a ({signal_1084, signal_775}), .c ({signal_1397, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_362 ( .s (signal_357), .b ({signal_877, signal_473}), .a ({signal_1087, signal_774}), .c ({signal_1398, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_363 ( .s (signal_357), .b ({signal_880, signal_472}), .a ({signal_1090, signal_773}), .c ({signal_1399, signal_777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_364 ( .s (signal_357), .b ({signal_883, signal_471}), .a ({signal_1093, signal_772}), .c ({signal_1400, signal_776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_373 ( .s (signal_357), .b ({signal_1305, signal_477}), .a ({signal_1096, signal_771}), .c ({signal_1401, signal_783}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_374 ( .s (signal_357), .b ({signal_1307, signal_476}), .a ({signal_1099, signal_770}), .c ({signal_1402, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_375 ( .s (signal_357), .b ({signal_1309, signal_475}), .a ({signal_1102, signal_769}), .c ({signal_1403, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_376 ( .s (signal_357), .b ({signal_1082, signal_695}), .a ({signal_1105, signal_768}), .c ({signal_1404, signal_780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_385 ( .s (signal_358), .b ({signal_1085, signal_694}), .a ({signal_1108, signal_767}), .c ({signal_1405, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_386 ( .s (signal_358), .b ({signal_1088, signal_693}), .a ({signal_1111, signal_766}), .c ({signal_1406, signal_786}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_387 ( .s (signal_358), .b ({signal_1091, signal_692}), .a ({signal_1114, signal_765}), .c ({signal_1407, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_388 ( .s (signal_358), .b ({signal_1094, signal_691}), .a ({signal_1117, signal_764}), .c ({signal_1408, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_397 ( .s (signal_358), .b ({signal_1097, signal_690}), .a ({signal_1120, signal_763}), .c ({signal_1409, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_398 ( .s (signal_358), .b ({signal_1100, signal_689}), .a ({signal_1123, signal_762}), .c ({signal_1410, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_399 ( .s (signal_358), .b ({signal_1103, signal_688}), .a ({signal_1126, signal_761}), .c ({signal_1411, signal_789}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_400 ( .s (signal_358), .b ({signal_1106, signal_687}), .a ({signal_1295, signal_760}), .c ({signal_1412, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_409 ( .s (signal_218), .b ({signal_1109, signal_686}), .a ({signal_1303, signal_759}), .c ({signal_1319, signal_795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_410 ( .s (signal_218), .b ({signal_1112, signal_685}), .a ({signal_1297, signal_758}), .c ({signal_1320, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_411 ( .s (signal_218), .b ({signal_1115, signal_684}), .a ({signal_1299, signal_757}), .c ({signal_1321, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_412 ( .s (signal_218), .b ({signal_1118, signal_683}), .a ({signal_1301, signal_756}), .c ({signal_1322, signal_792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_421 ( .s (signal_218), .b ({signal_1121, signal_682}), .a ({signal_1129, signal_755}), .c ({signal_1323, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_422 ( .s (signal_218), .b ({signal_1124, signal_681}), .a ({signal_1132, signal_754}), .c ({signal_1324, signal_798}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_423 ( .s (signal_218), .b ({signal_1080, signal_680}), .a ({signal_1135, signal_753}), .c ({signal_1325, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_424 ( .s (signal_218), .b ({signal_1292, signal_679}), .a ({signal_1138, signal_752}), .c ({signal_1326, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_433 ( .s (signal_357), .b ({signal_1078, signal_678}), .a ({signal_1141, signal_751}), .c ({signal_1413, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_434 ( .s (signal_357), .b ({signal_1076, signal_677}), .a ({signal_1144, signal_750}), .c ({signal_1414, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_435 ( .s (signal_357), .b ({signal_1074, signal_676}), .a ({signal_1147, signal_749}), .c ({signal_1415, signal_801}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_436 ( .s (signal_357), .b ({signal_1127, signal_675}), .a ({signal_1150, signal_748}), .c ({signal_1416, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_445 ( .s (signal_357), .b ({signal_1130, signal_674}), .a ({signal_1153, signal_747}), .c ({signal_1417, signal_807}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_446 ( .s (signal_357), .b ({signal_1133, signal_673}), .a ({signal_1156, signal_746}), .c ({signal_1418, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_447 ( .s (signal_357), .b ({signal_1136, signal_672}), .a ({signal_1159, signal_745}), .c ({signal_1419, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_448 ( .s (signal_357), .b ({signal_1139, signal_671}), .a ({signal_1162, signal_744}), .c ({signal_1420, signal_804}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_457 ( .s (signal_357), .b ({signal_1142, signal_670}), .a ({signal_1165, signal_743}), .c ({signal_1421, signal_811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_458 ( .s (signal_357), .b ({signal_1145, signal_669}), .a ({signal_1168, signal_742}), .c ({signal_1422, signal_810}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_459 ( .s (signal_357), .b ({signal_1148, signal_668}), .a ({signal_1171, signal_741}), .c ({signal_1423, signal_809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_460 ( .s (signal_357), .b ({signal_1151, signal_667}), .a ({signal_1174, signal_740}), .c ({signal_1424, signal_808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_469 ( .s (signal_357), .b ({signal_1154, signal_666}), .a ({signal_1177, signal_739}), .c ({signal_1425, signal_815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_470 ( .s (signal_357), .b ({signal_1157, signal_665}), .a ({signal_1180, signal_738}), .c ({signal_1426, signal_814}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_471 ( .s (signal_357), .b ({signal_1160, signal_664}), .a ({signal_1183, signal_737}), .c ({signal_1427, signal_813}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_472 ( .s (signal_357), .b ({signal_1163, signal_663}), .a ({signal_1186, signal_736}), .c ({signal_1428, signal_812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_481 ( .s (signal_357), .b ({signal_1166, signal_662}), .a ({signal_1189, signal_735}), .c ({signal_1429, signal_819}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_482 ( .s (signal_357), .b ({signal_1169, signal_661}), .a ({signal_1192, signal_734}), .c ({signal_1430, signal_818}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_483 ( .s (signal_357), .b ({signal_1172, signal_660}), .a ({signal_1195, signal_733}), .c ({signal_1431, signal_817}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_484 ( .s (signal_357), .b ({signal_1175, signal_659}), .a ({signal_1198, signal_732}), .c ({signal_1432, signal_816}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_493 ( .s (signal_357), .b ({signal_1178, signal_658}), .a ({signal_1201, signal_731}), .c ({signal_1433, signal_823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_494 ( .s (signal_357), .b ({signal_1181, signal_657}), .a ({signal_1204, signal_730}), .c ({signal_1434, signal_822}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_495 ( .s (signal_357), .b ({signal_1184, signal_656}), .a ({signal_1207, signal_729}), .c ({signal_1435, signal_821}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_496 ( .s (signal_357), .b ({signal_1187, signal_655}), .a ({signal_1210, signal_728}), .c ({signal_1436, signal_820}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_505 ( .s (signal_357), .b ({signal_1190, signal_654}), .a ({signal_1213, signal_727}), .c ({signal_1437, signal_827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_506 ( .s (signal_357), .b ({signal_1193, signal_653}), .a ({signal_1216, signal_726}), .c ({signal_1438, signal_826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_507 ( .s (signal_357), .b ({signal_1196, signal_652}), .a ({signal_1219, signal_725}), .c ({signal_1439, signal_825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_508 ( .s (signal_357), .b ({signal_1199, signal_651}), .a ({signal_1222, signal_724}), .c ({signal_1440, signal_824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_517 ( .s (signal_358), .b ({signal_1202, signal_650}), .a ({signal_1225, signal_723}), .c ({signal_1441, signal_831}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_518 ( .s (signal_358), .b ({signal_1205, signal_649}), .a ({signal_1228, signal_722}), .c ({signal_1442, signal_830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_519 ( .s (signal_358), .b ({signal_1208, signal_648}), .a ({signal_1231, signal_721}), .c ({signal_1443, signal_829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_520 ( .s (signal_358), .b ({signal_1211, signal_647}), .a ({signal_1234, signal_720}), .c ({signal_1444, signal_828}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_529 ( .s (signal_358), .b ({signal_1214, signal_646}), .a ({signal_1237, signal_719}), .c ({signal_1445, signal_835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_530 ( .s (signal_358), .b ({signal_1217, signal_645}), .a ({signal_1240, signal_718}), .c ({signal_1446, signal_834}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_531 ( .s (signal_358), .b ({signal_1220, signal_644}), .a ({signal_1243, signal_717}), .c ({signal_1447, signal_833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_532 ( .s (signal_358), .b ({signal_1223, signal_643}), .a ({signal_1246, signal_716}), .c ({signal_1448, signal_832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_541 ( .s (signal_358), .b ({signal_1226, signal_642}), .a ({signal_1249, signal_715}), .c ({signal_1449, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_542 ( .s (signal_358), .b ({signal_1229, signal_641}), .a ({signal_1252, signal_714}), .c ({signal_1450, signal_838}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_543 ( .s (signal_358), .b ({signal_1232, signal_640}), .a ({signal_1255, signal_713}), .c ({signal_1451, signal_837}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_544 ( .s (signal_358), .b ({signal_1235, signal_639}), .a ({signal_1258, signal_712}), .c ({signal_1452, signal_836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_553 ( .s (signal_358), .b ({signal_1238, signal_638}), .a ({signal_1261, signal_711}), .c ({signal_1453, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_554 ( .s (signal_358), .b ({signal_1241, signal_637}), .a ({signal_1264, signal_710}), .c ({signal_1454, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_555 ( .s (signal_358), .b ({signal_1244, signal_636}), .a ({signal_1267, signal_709}), .c ({signal_1455, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_556 ( .s (signal_358), .b ({signal_1247, signal_635}), .a ({signal_1270, signal_708}), .c ({signal_1456, signal_840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_565 ( .s (signal_358), .b ({signal_1250, signal_634}), .a ({signal_1273, signal_707}), .c ({signal_1457, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_566 ( .s (signal_358), .b ({signal_1253, signal_633}), .a ({signal_1276, signal_706}), .c ({signal_1458, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_567 ( .s (signal_358), .b ({signal_1256, signal_632}), .a ({signal_1279, signal_705}), .c ({signal_1459, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_568 ( .s (signal_358), .b ({signal_1259, signal_631}), .a ({signal_1282, signal_704}), .c ({signal_1460, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_577 ( .s (signal_358), .b ({signal_1262, signal_630}), .a ({signal_1285, signal_703}), .c ({signal_1461, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_578 ( .s (signal_358), .b ({signal_1265, signal_629}), .a ({signal_1287, signal_702}), .c ({signal_1462, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_579 ( .s (signal_358), .b ({signal_1268, signal_628}), .a ({signal_1289, signal_701}), .c ({signal_1463, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_580 ( .s (signal_358), .b ({signal_1271, signal_627}), .a ({signal_1291, signal_700}), .c ({signal_1464, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_593 ( .s (reset), .b ({signal_1082, signal_695}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1084, signal_775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_594 ( .s (reset), .b ({signal_1085, signal_694}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1087, signal_774}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_595 ( .s (reset), .b ({signal_1088, signal_693}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1090, signal_773}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_596 ( .s (reset), .b ({signal_1091, signal_692}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1093, signal_772}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_597 ( .s (reset), .b ({signal_1094, signal_691}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1096, signal_771}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_598 ( .s (reset), .b ({signal_1097, signal_690}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1099, signal_770}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_599 ( .s (reset), .b ({signal_1100, signal_689}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1102, signal_769}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_600 ( .s (reset), .b ({signal_1103, signal_688}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1105, signal_768}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_601 ( .s (reset), .b ({signal_1106, signal_687}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1108, signal_767}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_602 ( .s (reset), .b ({signal_1109, signal_686}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1111, signal_766}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_603 ( .s (reset), .b ({signal_1112, signal_685}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1114, signal_765}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_604 ( .s (reset), .b ({signal_1115, signal_684}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1117, signal_764}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_605 ( .s (reset), .b ({signal_1118, signal_683}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1120, signal_763}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_606 ( .s (reset), .b ({signal_1121, signal_682}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1123, signal_762}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_607 ( .s (reset), .b ({signal_1124, signal_681}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1126, signal_761}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_608 ( .s (reset), .b ({signal_1081, signal_622}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1295, signal_760}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_609 ( .s (reset), .b ({signal_1293, signal_621}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1303, signal_759}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_610 ( .s (reset), .b ({signal_1079, signal_620}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1297, signal_758}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_611 ( .s (reset), .b ({signal_1077, signal_619}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1299, signal_757}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_612 ( .s (reset), .b ({signal_1075, signal_618}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1301, signal_756}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_613 ( .s (reset), .b ({signal_1127, signal_675}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1129, signal_755}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_614 ( .s (reset), .b ({signal_1130, signal_674}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1132, signal_754}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_615 ( .s (reset), .b ({signal_1133, signal_673}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1135, signal_753}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_616 ( .s (reset), .b ({signal_1136, signal_672}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1138, signal_752}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_617 ( .s (reset), .b ({signal_1139, signal_671}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1141, signal_751}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_618 ( .s (reset), .b ({signal_1142, signal_670}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1144, signal_750}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_619 ( .s (reset), .b ({signal_1145, signal_669}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1147, signal_749}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_620 ( .s (reset), .b ({signal_1148, signal_668}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1150, signal_748}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_621 ( .s (reset), .b ({signal_1151, signal_667}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1153, signal_747}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_622 ( .s (reset), .b ({signal_1154, signal_666}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1156, signal_746}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_623 ( .s (reset), .b ({signal_1157, signal_665}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1159, signal_745}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_624 ( .s (reset), .b ({signal_1160, signal_664}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1162, signal_744}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_625 ( .s (reset), .b ({signal_1163, signal_663}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1165, signal_743}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_626 ( .s (reset), .b ({signal_1166, signal_662}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1168, signal_742}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_627 ( .s (reset), .b ({signal_1169, signal_661}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1171, signal_741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_628 ( .s (reset), .b ({signal_1172, signal_660}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1174, signal_740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_629 ( .s (reset), .b ({signal_1175, signal_659}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1177, signal_739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_630 ( .s (reset), .b ({signal_1178, signal_658}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1180, signal_738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_631 ( .s (reset), .b ({signal_1181, signal_657}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1183, signal_737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_632 ( .s (reset), .b ({signal_1184, signal_656}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1186, signal_736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_633 ( .s (reset), .b ({signal_1187, signal_655}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1189, signal_735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_634 ( .s (reset), .b ({signal_1190, signal_654}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1192, signal_734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_635 ( .s (reset), .b ({signal_1193, signal_653}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1195, signal_733}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_636 ( .s (reset), .b ({signal_1196, signal_652}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1198, signal_732}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_637 ( .s (reset), .b ({signal_1199, signal_651}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1201, signal_731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_638 ( .s (reset), .b ({signal_1202, signal_650}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1204, signal_730}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_639 ( .s (reset), .b ({signal_1205, signal_649}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1207, signal_729}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_640 ( .s (reset), .b ({signal_1208, signal_648}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1210, signal_728}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_641 ( .s (reset), .b ({signal_1211, signal_647}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1213, signal_727}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_642 ( .s (reset), .b ({signal_1214, signal_646}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1216, signal_726}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_643 ( .s (reset), .b ({signal_1217, signal_645}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1219, signal_725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_644 ( .s (reset), .b ({signal_1220, signal_644}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1222, signal_724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_645 ( .s (reset), .b ({signal_1223, signal_643}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1225, signal_723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_646 ( .s (reset), .b ({signal_1226, signal_642}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1228, signal_722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_647 ( .s (reset), .b ({signal_1229, signal_641}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1231, signal_721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_648 ( .s (reset), .b ({signal_1232, signal_640}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1234, signal_720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_649 ( .s (reset), .b ({signal_1235, signal_639}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1237, signal_719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_650 ( .s (reset), .b ({signal_1238, signal_638}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1240, signal_718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_651 ( .s (reset), .b ({signal_1241, signal_637}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1243, signal_717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_652 ( .s (reset), .b ({signal_1244, signal_636}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1246, signal_716}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_653 ( .s (reset), .b ({signal_1247, signal_635}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1249, signal_715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_654 ( .s (reset), .b ({signal_1250, signal_634}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1252, signal_714}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_655 ( .s (reset), .b ({signal_1253, signal_633}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1255, signal_713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_656 ( .s (reset), .b ({signal_1256, signal_632}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1258, signal_712}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_657 ( .s (reset), .b ({signal_1259, signal_631}), .a ({key_s1[64], key_s0[64]}), .c ({signal_1261, signal_711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_658 ( .s (reset), .b ({signal_1262, signal_630}), .a ({key_s1[65], key_s0[65]}), .c ({signal_1264, signal_710}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_659 ( .s (reset), .b ({signal_1265, signal_629}), .a ({key_s1[66], key_s0[66]}), .c ({signal_1267, signal_709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_660 ( .s (reset), .b ({signal_1268, signal_628}), .a ({key_s1[67], key_s0[67]}), .c ({signal_1270, signal_708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_661 ( .s (reset), .b ({signal_1271, signal_627}), .a ({key_s1[68], key_s0[68]}), .c ({signal_1273, signal_707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_662 ( .s (reset), .b ({signal_1274, signal_626}), .a ({key_s1[69], key_s0[69]}), .c ({signal_1276, signal_706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_663 ( .s (reset), .b ({signal_1277, signal_625}), .a ({key_s1[70], key_s0[70]}), .c ({signal_1279, signal_705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_664 ( .s (reset), .b ({signal_1280, signal_624}), .a ({key_s1[71], key_s0[71]}), .c ({signal_1282, signal_704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_665 ( .s (reset), .b ({signal_1283, signal_623}), .a ({key_s1[72], key_s0[72]}), .c ({signal_1285, signal_703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_666 ( .s (reset), .b ({signal_874, signal_474}), .a ({key_s1[73], key_s0[73]}), .c ({signal_1287, signal_702}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_667 ( .s (reset), .b ({signal_877, signal_473}), .a ({key_s1[74], key_s0[74]}), .c ({signal_1289, signal_701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_668 ( .s (reset), .b ({signal_880, signal_472}), .a ({key_s1[75], key_s0[75]}), .c ({signal_1291, signal_700}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_696 ( .s (signal_217), .b ({signal_876, signal_485}), .a ({signal_883, signal_471}), .c ({signal_1304, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_697 ( .s (signal_217), .b ({signal_879, signal_484}), .a ({signal_1305, signal_477}), .c ({signal_1306, signal_480}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_698 ( .s (signal_217), .b ({signal_882, signal_483}), .a ({signal_1307, signal_476}), .c ({signal_1308, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_699 ( .s (signal_217), .b ({signal_885, signal_482}), .a ({signal_1309, signal_475}), .c ({signal_1310, signal_478}) ) ;
    ClockGatingController #(9) cell_726 ( .clk (clk), .rst (reset), .GatedClk (signal_1512), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_704 ( .s ({signal_1306, signal_480}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[0]), .c ({signal_1311, signal_856}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_705 ( .s ({signal_1308, signal_479}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[1]), .c ({signal_1312, signal_857}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_706 ( .s ({signal_1308, signal_479}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[2]), .c ({signal_1313, signal_858}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_707 ( .s ({signal_1306, signal_480}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[3]), .c ({signal_1314, signal_859}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_708 ( .s ({signal_1310, signal_478}), .b ({signal_1314, signal_859}), .a ({signal_1313, signal_858}), .clk (clk), .r (Fresh[4]), .c ({signal_1327, signal_860}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_709 ( .s ({signal_1308, signal_479}), .b ({signal_1314, signal_859}), .a ({signal_1311, signal_856}), .clk (clk), .r (Fresh[5]), .c ({signal_1328, signal_861}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_710 ( .s ({signal_1308, signal_479}), .b ({signal_1311, signal_856}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[6]), .c ({signal_1329, signal_862}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_711 ( .s ({signal_1308, signal_479}), .b ({signal_1314, signal_859}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[7]), .c ({signal_1330, signal_863}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_712 ( .s ({signal_1308, signal_479}), .b ({1'b0, 1'b0}), .a ({signal_1314, signal_859}), .clk (clk), .r (Fresh[8]), .c ({signal_1331, signal_864}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_713 ( .s ({signal_1310, signal_478}), .b ({signal_1311, signal_856}), .a ({signal_1312, signal_857}), .clk (clk), .r (Fresh[9]), .c ({signal_1332, signal_865}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_714 ( .s ({signal_1308, signal_479}), .b ({1'b0, 1'b1}), .a ({signal_1311, signal_856}), .clk (clk), .r (Fresh[10]), .c ({signal_1333, signal_866}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_715 ( .s ({signal_1308, signal_479}), .b ({signal_1311, signal_856}), .a ({signal_1314, signal_859}), .clk (clk), .r (Fresh[11]), .c ({signal_1334, signal_867}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_716 ( .s ({signal_1310, signal_478}), .b ({signal_1312, signal_857}), .a ({signal_1334, signal_867}), .clk (clk), .r (Fresh[12]), .c ({signal_1335, signal_868}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_717 ( .s ({signal_1310, signal_478}), .b ({signal_1331, signal_864}), .a ({signal_1333, signal_866}), .clk (clk), .r (Fresh[13]), .c ({signal_1336, signal_869}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_718 ( .s ({signal_1310, signal_478}), .b ({signal_1333, signal_866}), .a ({signal_1331, signal_864}), .clk (clk), .r (Fresh[14]), .c ({signal_1337, signal_870}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_719 ( .s ({signal_1310, signal_478}), .b ({signal_1329, signal_862}), .a ({signal_1330, signal_863}), .clk (clk), .r (Fresh[15]), .c ({signal_1338, signal_871}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_720 ( .s ({signal_1310, signal_478}), .b ({signal_1330, signal_863}), .a ({signal_1329, signal_862}), .clk (clk), .r (Fresh[16]), .c ({signal_1339, signal_872}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_721 ( .s ({signal_1310, signal_478}), .b ({signal_1328, signal_861}), .a ({signal_1314, signal_859}), .clk (clk), .r (Fresh[17]), .c ({signal_1340, signal_873}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_89 ( .s (signal_218), .b ({signal_1476, signal_466}), .a ({signal_888, signal_553}), .c ({signal_1479, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_90 ( .s (signal_218), .b ({signal_1477, signal_465}), .a ({signal_891, signal_552}), .c ({signal_1480, signal_556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_91 ( .s (signal_218), .b ({signal_1478, signal_464}), .a ({signal_894, signal_551}), .c ({signal_1481, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_92 ( .s (signal_218), .b ({signal_1487, signal_463}), .a ({signal_897, signal_550}), .c ({signal_1488, signal_554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_589 ( .s (signal_358), .b ({signal_1274, signal_626}), .a ({signal_1470, signal_699}), .c ({signal_1482, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_590 ( .s (signal_358), .b ({signal_1277, signal_625}), .a ({signal_1472, signal_698}), .c ({signal_1483, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_591 ( .s (signal_358), .b ({signal_1280, signal_624}), .a ({signal_1474, signal_697}), .c ({signal_1484, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_592 ( .s (signal_358), .b ({signal_1283, signal_623}), .a ({signal_1486, signal_696}), .c ({signal_1489, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_669 ( .s (reset), .b ({signal_1467, signal_470}), .a ({key_s1[76], key_s0[76]}), .c ({signal_1470, signal_699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_670 ( .s (reset), .b ({signal_1466, signal_469}), .a ({key_s1[77], key_s0[77]}), .c ({signal_1472, signal_698}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_671 ( .s (reset), .b ({signal_1465, signal_468}), .a ({key_s1[78], key_s0[78]}), .c ({signal_1474, signal_697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_672 ( .s (reset), .b ({signal_1475, signal_467}), .a ({key_s1[79], key_s0[79]}), .c ({signal_1486, signal_696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_691 ( .a ({signal_1304, signal_481}), .b ({signal_1468, signal_443}), .c ({signal_1475, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_700 ( .s (signal_219), .b ({signal_1467, signal_470}), .a ({signal_876, signal_485}), .c ({signal_1476, signal_466}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_701 ( .s (signal_219), .b ({signal_1466, signal_469}), .a ({signal_879, signal_484}), .c ({signal_1477, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_702 ( .s (signal_219), .b ({signal_1465, signal_468}), .a ({signal_882, signal_483}), .c ({signal_1478, signal_464}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_703 ( .s (signal_219), .b ({signal_1475, signal_467}), .a ({signal_885, signal_482}), .c ({signal_1487, signal_463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_722 ( .s ({signal_1304, signal_481}), .b ({signal_1335, signal_868}), .a ({signal_1340, signal_873}), .clk (clk), .r (Fresh[18]), .c ({signal_1465, signal_468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_723 ( .s ({signal_1304, signal_481}), .b ({signal_1332, signal_865}), .a ({signal_1338, signal_871}), .clk (clk), .r (Fresh[19]), .c ({signal_1466, signal_469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_724 ( .s ({signal_1304, signal_481}), .b ({signal_1336, signal_869}), .a ({signal_1337, signal_870}), .clk (clk), .r (Fresh[20]), .c ({signal_1467, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_725 ( .s ({signal_1304, signal_481}), .b ({signal_1339, signal_872}), .a ({signal_1327, signal_860}), .clk (clk), .r (Fresh[21]), .c ({signal_1468, signal_443}) ) ;

    /* register cells */
    DFF_X1 cell_53 ( .CK (signal_1512), .D (signal_271), .Q (signal_458), .QN () ) ;
    DFF_X1 cell_55 ( .CK (signal_1512), .D (signal_270), .Q (signal_460), .QN () ) ;
    DFF_X1 cell_57 ( .CK (signal_1512), .D (signal_269), .Q (signal_462), .QN () ) ;
    DFF_X1 cell_59 ( .CK (signal_1512), .D (signal_268), .Q (signal_459), .QN () ) ;
    DFF_X1 cell_61 ( .CK (signal_1512), .D (signal_266), .Q (signal_265), .QN () ) ;
    DFF_X1 cell_75 ( .CK (signal_1512), .D (signal_285), .Q (signal_487), .QN () ) ;
    DFF_X1 cell_77 ( .CK (signal_1512), .D (signal_284), .Q (signal_489), .QN () ) ;
    DFF_X1 cell_79 ( .CK (signal_1512), .D (signal_283), .Q (signal_486), .QN () ) ;
    DFF_X1 cell_81 ( .CK (signal_1512), .D (signal_282), .Q (signal_488), .QN () ) ;
    DFF_X1 cell_83 ( .CK (signal_1512), .D (signal_236), .Q (signal_234), .QN () ) ;
    DFF_X1 cell_85 ( .CK (signal_1512), .D (signal_233), .Q (signal_235), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_94 ( .clk (signal_1512), .D ({signal_1479, signal_557}), .Q ({data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_96 ( .clk (signal_1512), .D ({signal_1481, signal_555}), .Q ({data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_98 ( .clk (signal_1512), .D ({signal_1480, signal_556}), .Q ({data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_100 ( .clk (signal_1512), .D ({signal_1488, signal_554}), .Q ({data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_102 ( .clk (signal_1512), .D ({signal_1318, signal_558}), .Q ({data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_104 ( .clk (signal_1512), .D ({signal_1317, signal_559}), .Q ({data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_106 ( .clk (signal_1512), .D ({signal_1316, signal_560}), .Q ({data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_108 ( .clk (signal_1512), .D ({signal_1315, signal_561}), .Q ({data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_114 ( .clk (signal_1512), .D ({signal_1344, signal_562}), .Q ({data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_116 ( .clk (signal_1512), .D ({signal_1343, signal_563}), .Q ({data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_118 ( .clk (signal_1512), .D ({signal_1342, signal_564}), .Q ({data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_120 ( .clk (signal_1512), .D ({signal_1341, signal_565}), .Q ({data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_126 ( .clk (signal_1512), .D ({signal_1348, signal_566}), .Q ({data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_128 ( .clk (signal_1512), .D ({signal_1347, signal_567}), .Q ({data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_130 ( .clk (signal_1512), .D ({signal_1346, signal_568}), .Q ({data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_132 ( .clk (signal_1512), .D ({signal_1345, signal_569}), .Q ({data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_138 ( .clk (signal_1512), .D ({signal_1352, signal_570}), .Q ({data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_140 ( .clk (signal_1512), .D ({signal_1351, signal_571}), .Q ({data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_142 ( .clk (signal_1512), .D ({signal_1350, signal_572}), .Q ({data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_144 ( .clk (signal_1512), .D ({signal_1349, signal_573}), .Q ({data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_150 ( .clk (signal_1512), .D ({signal_1356, signal_574}), .Q ({data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_152 ( .clk (signal_1512), .D ({signal_1355, signal_575}), .Q ({data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_154 ( .clk (signal_1512), .D ({signal_1354, signal_576}), .Q ({data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_156 ( .clk (signal_1512), .D ({signal_1353, signal_577}), .Q ({data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_162 ( .clk (signal_1512), .D ({signal_1360, signal_578}), .Q ({data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_164 ( .clk (signal_1512), .D ({signal_1359, signal_579}), .Q ({data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_166 ( .clk (signal_1512), .D ({signal_1358, signal_580}), .Q ({data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_168 ( .clk (signal_1512), .D ({signal_1357, signal_581}), .Q ({data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_174 ( .clk (signal_1512), .D ({signal_1364, signal_582}), .Q ({data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_176 ( .clk (signal_1512), .D ({signal_1363, signal_583}), .Q ({data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_178 ( .clk (signal_1512), .D ({signal_1362, signal_584}), .Q ({data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_180 ( .clk (signal_1512), .D ({signal_1361, signal_585}), .Q ({data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_186 ( .clk (signal_1512), .D ({signal_1368, signal_586}), .Q ({data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_188 ( .clk (signal_1512), .D ({signal_1367, signal_587}), .Q ({data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_190 ( .clk (signal_1512), .D ({signal_1366, signal_588}), .Q ({data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_192 ( .clk (signal_1512), .D ({signal_1365, signal_589}), .Q ({data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_198 ( .clk (signal_1512), .D ({signal_1372, signal_590}), .Q ({data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_200 ( .clk (signal_1512), .D ({signal_1371, signal_591}), .Q ({data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_202 ( .clk (signal_1512), .D ({signal_1370, signal_592}), .Q ({data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_204 ( .clk (signal_1512), .D ({signal_1369, signal_593}), .Q ({data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_210 ( .clk (signal_1512), .D ({signal_1376, signal_594}), .Q ({data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_212 ( .clk (signal_1512), .D ({signal_1375, signal_595}), .Q ({data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_214 ( .clk (signal_1512), .D ({signal_1374, signal_596}), .Q ({data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_216 ( .clk (signal_1512), .D ({signal_1373, signal_597}), .Q ({data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_222 ( .clk (signal_1512), .D ({signal_1380, signal_598}), .Q ({data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_224 ( .clk (signal_1512), .D ({signal_1379, signal_599}), .Q ({data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_226 ( .clk (signal_1512), .D ({signal_1378, signal_600}), .Q ({data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_228 ( .clk (signal_1512), .D ({signal_1377, signal_601}), .Q ({data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_234 ( .clk (signal_1512), .D ({signal_1384, signal_602}), .Q ({data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_236 ( .clk (signal_1512), .D ({signal_1383, signal_603}), .Q ({data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_238 ( .clk (signal_1512), .D ({signal_1382, signal_604}), .Q ({data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_240 ( .clk (signal_1512), .D ({signal_1381, signal_605}), .Q ({data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_246 ( .clk (signal_1512), .D ({signal_1388, signal_606}), .Q ({data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_248 ( .clk (signal_1512), .D ({signal_1387, signal_607}), .Q ({data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_250 ( .clk (signal_1512), .D ({signal_1386, signal_608}), .Q ({data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_252 ( .clk (signal_1512), .D ({signal_1385, signal_609}), .Q ({data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_258 ( .clk (signal_1512), .D ({signal_1392, signal_610}), .Q ({data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_260 ( .clk (signal_1512), .D ({signal_1391, signal_611}), .Q ({data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_262 ( .clk (signal_1512), .D ({signal_1390, signal_612}), .Q ({data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_264 ( .clk (signal_1512), .D ({signal_1389, signal_613}), .Q ({data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_270 ( .clk (signal_1512), .D ({signal_1396, signal_614}), .Q ({data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_272 ( .clk (signal_1512), .D ({signal_1395, signal_615}), .Q ({data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_274 ( .clk (signal_1512), .D ({signal_1394, signal_616}), .Q ({data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_276 ( .clk (signal_1512), .D ({signal_1393, signal_617}), .Q ({data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_354 ( .clk (signal_1512), .D ({signal_1400, signal_776}), .Q ({signal_1082, signal_695}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_356 ( .clk (signal_1512), .D ({signal_1399, signal_777}), .Q ({signal_1309, signal_475}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_358 ( .clk (signal_1512), .D ({signal_1398, signal_778}), .Q ({signal_1307, signal_476}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_360 ( .clk (signal_1512), .D ({signal_1397, signal_779}), .Q ({signal_1305, signal_477}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_366 ( .clk (signal_1512), .D ({signal_1404, signal_780}), .Q ({signal_1094, signal_691}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_368 ( .clk (signal_1512), .D ({signal_1403, signal_781}), .Q ({signal_1091, signal_692}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_370 ( .clk (signal_1512), .D ({signal_1402, signal_782}), .Q ({signal_1088, signal_693}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_372 ( .clk (signal_1512), .D ({signal_1401, signal_783}), .Q ({signal_1085, signal_694}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_378 ( .clk (signal_1512), .D ({signal_1408, signal_784}), .Q ({signal_1106, signal_687}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_380 ( .clk (signal_1512), .D ({signal_1407, signal_785}), .Q ({signal_1103, signal_688}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_382 ( .clk (signal_1512), .D ({signal_1406, signal_786}), .Q ({signal_1100, signal_689}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_384 ( .clk (signal_1512), .D ({signal_1405, signal_787}), .Q ({signal_1097, signal_690}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_390 ( .clk (signal_1512), .D ({signal_1412, signal_788}), .Q ({signal_1118, signal_683}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_392 ( .clk (signal_1512), .D ({signal_1411, signal_789}), .Q ({signal_1115, signal_684}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_394 ( .clk (signal_1512), .D ({signal_1410, signal_790}), .Q ({signal_1112, signal_685}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_396 ( .clk (signal_1512), .D ({signal_1409, signal_791}), .Q ({signal_1109, signal_686}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_402 ( .clk (signal_1512), .D ({signal_1322, signal_792}), .Q ({signal_1292, signal_679}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_404 ( .clk (signal_1512), .D ({signal_1321, signal_793}), .Q ({signal_1080, signal_680}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_406 ( .clk (signal_1512), .D ({signal_1320, signal_794}), .Q ({signal_1124, signal_681}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_408 ( .clk (signal_1512), .D ({signal_1319, signal_795}), .Q ({signal_1121, signal_682}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_414 ( .clk (signal_1512), .D ({signal_1326, signal_796}), .Q ({signal_1127, signal_675}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_416 ( .clk (signal_1512), .D ({signal_1325, signal_797}), .Q ({signal_1074, signal_676}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_418 ( .clk (signal_1512), .D ({signal_1324, signal_798}), .Q ({signal_1076, signal_677}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_420 ( .clk (signal_1512), .D ({signal_1323, signal_799}), .Q ({signal_1078, signal_678}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_426 ( .clk (signal_1512), .D ({signal_1416, signal_800}), .Q ({signal_1139, signal_671}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_428 ( .clk (signal_1512), .D ({signal_1415, signal_801}), .Q ({signal_1136, signal_672}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_430 ( .clk (signal_1512), .D ({signal_1414, signal_802}), .Q ({signal_1133, signal_673}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_432 ( .clk (signal_1512), .D ({signal_1413, signal_803}), .Q ({signal_1130, signal_674}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_438 ( .clk (signal_1512), .D ({signal_1420, signal_804}), .Q ({signal_1151, signal_667}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_440 ( .clk (signal_1512), .D ({signal_1419, signal_805}), .Q ({signal_1148, signal_668}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_442 ( .clk (signal_1512), .D ({signal_1418, signal_806}), .Q ({signal_1145, signal_669}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_444 ( .clk (signal_1512), .D ({signal_1417, signal_807}), .Q ({signal_1142, signal_670}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_450 ( .clk (signal_1512), .D ({signal_1424, signal_808}), .Q ({signal_1163, signal_663}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_452 ( .clk (signal_1512), .D ({signal_1423, signal_809}), .Q ({signal_1160, signal_664}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_454 ( .clk (signal_1512), .D ({signal_1422, signal_810}), .Q ({signal_1157, signal_665}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_456 ( .clk (signal_1512), .D ({signal_1421, signal_811}), .Q ({signal_1154, signal_666}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_462 ( .clk (signal_1512), .D ({signal_1428, signal_812}), .Q ({signal_1175, signal_659}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_464 ( .clk (signal_1512), .D ({signal_1427, signal_813}), .Q ({signal_1172, signal_660}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_466 ( .clk (signal_1512), .D ({signal_1426, signal_814}), .Q ({signal_1169, signal_661}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_468 ( .clk (signal_1512), .D ({signal_1425, signal_815}), .Q ({signal_1166, signal_662}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_474 ( .clk (signal_1512), .D ({signal_1432, signal_816}), .Q ({signal_1187, signal_655}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_476 ( .clk (signal_1512), .D ({signal_1431, signal_817}), .Q ({signal_1184, signal_656}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_478 ( .clk (signal_1512), .D ({signal_1430, signal_818}), .Q ({signal_1181, signal_657}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_480 ( .clk (signal_1512), .D ({signal_1429, signal_819}), .Q ({signal_1178, signal_658}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_486 ( .clk (signal_1512), .D ({signal_1436, signal_820}), .Q ({signal_1199, signal_651}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_488 ( .clk (signal_1512), .D ({signal_1435, signal_821}), .Q ({signal_1196, signal_652}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_490 ( .clk (signal_1512), .D ({signal_1434, signal_822}), .Q ({signal_1193, signal_653}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_492 ( .clk (signal_1512), .D ({signal_1433, signal_823}), .Q ({signal_1190, signal_654}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_498 ( .clk (signal_1512), .D ({signal_1440, signal_824}), .Q ({signal_1211, signal_647}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_500 ( .clk (signal_1512), .D ({signal_1439, signal_825}), .Q ({signal_1208, signal_648}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_502 ( .clk (signal_1512), .D ({signal_1438, signal_826}), .Q ({signal_1205, signal_649}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_504 ( .clk (signal_1512), .D ({signal_1437, signal_827}), .Q ({signal_1202, signal_650}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_510 ( .clk (signal_1512), .D ({signal_1444, signal_828}), .Q ({signal_1223, signal_643}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_512 ( .clk (signal_1512), .D ({signal_1443, signal_829}), .Q ({signal_1220, signal_644}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_514 ( .clk (signal_1512), .D ({signal_1442, signal_830}), .Q ({signal_1217, signal_645}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_516 ( .clk (signal_1512), .D ({signal_1441, signal_831}), .Q ({signal_1214, signal_646}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_522 ( .clk (signal_1512), .D ({signal_1448, signal_832}), .Q ({signal_1235, signal_639}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_524 ( .clk (signal_1512), .D ({signal_1447, signal_833}), .Q ({signal_1232, signal_640}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_526 ( .clk (signal_1512), .D ({signal_1446, signal_834}), .Q ({signal_1229, signal_641}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_528 ( .clk (signal_1512), .D ({signal_1445, signal_835}), .Q ({signal_1226, signal_642}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_534 ( .clk (signal_1512), .D ({signal_1452, signal_836}), .Q ({signal_1247, signal_635}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_536 ( .clk (signal_1512), .D ({signal_1451, signal_837}), .Q ({signal_1244, signal_636}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_538 ( .clk (signal_1512), .D ({signal_1450, signal_838}), .Q ({signal_1241, signal_637}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_540 ( .clk (signal_1512), .D ({signal_1449, signal_839}), .Q ({signal_1238, signal_638}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_546 ( .clk (signal_1512), .D ({signal_1456, signal_840}), .Q ({signal_1259, signal_631}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_548 ( .clk (signal_1512), .D ({signal_1455, signal_841}), .Q ({signal_1256, signal_632}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_550 ( .clk (signal_1512), .D ({signal_1454, signal_842}), .Q ({signal_1253, signal_633}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_552 ( .clk (signal_1512), .D ({signal_1453, signal_843}), .Q ({signal_1250, signal_634}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_558 ( .clk (signal_1512), .D ({signal_1460, signal_844}), .Q ({signal_1271, signal_627}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_560 ( .clk (signal_1512), .D ({signal_1459, signal_845}), .Q ({signal_1268, signal_628}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_562 ( .clk (signal_1512), .D ({signal_1458, signal_846}), .Q ({signal_1265, signal_629}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_564 ( .clk (signal_1512), .D ({signal_1457, signal_847}), .Q ({signal_1262, signal_630}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_570 ( .clk (signal_1512), .D ({signal_1464, signal_848}), .Q ({signal_1283, signal_623}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_572 ( .clk (signal_1512), .D ({signal_1463, signal_849}), .Q ({signal_1280, signal_624}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_574 ( .clk (signal_1512), .D ({signal_1462, signal_850}), .Q ({signal_1277, signal_625}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_576 ( .clk (signal_1512), .D ({signal_1461, signal_851}), .Q ({signal_1274, signal_626}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_582 ( .clk (signal_1512), .D ({signal_1489, signal_852}), .Q ({signal_883, signal_471}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_584 ( .clk (signal_1512), .D ({signal_1484, signal_853}), .Q ({signal_880, signal_472}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_586 ( .clk (signal_1512), .D ({signal_1483, signal_854}), .Q ({signal_877, signal_473}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_588 ( .clk (signal_1512), .D ({signal_1482, signal_855}), .Q ({signal_874, signal_474}) ) ;
endmodule
