/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [3:0] X_s3 ;
    input [23:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    output [3:0] Y_s3 ;
    wire Q0 ;
    wire Q1 ;
    wire T0 ;
    wire Q2 ;
    wire T1 ;
    wire Q4 ;
    wire T2 ;
    wire L0 ;
    wire Q6 ;
    wire L1 ;
    wire Q7 ;
    wire T3 ;
    wire L2 ;
    wire L2_T1 ;
    wire L3 ;
    wire n2 ;
    wire [2:1] XX ;
    wire [3:0] YY ;
    wire new_AGEMA_signal_40 ;
    wire new_AGEMA_signal_41 ;
    wire new_AGEMA_signal_42 ;
    wire new_AGEMA_signal_46 ;
    wire new_AGEMA_signal_47 ;
    wire new_AGEMA_signal_48 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_53 ;
    wire new_AGEMA_signal_54 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_61 ;
    wire new_AGEMA_signal_62 ;
    wire new_AGEMA_signal_63 ;
    wire new_AGEMA_signal_64 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_89 ;
    wire new_AGEMA_signal_90 ;
    wire new_AGEMA_signal_91 ;
    wire new_AGEMA_signal_92 ;
    wire new_AGEMA_signal_93 ;
    wire new_AGEMA_signal_94 ;
    wire new_AGEMA_signal_95 ;
    wire new_AGEMA_signal_96 ;
    wire new_AGEMA_signal_97 ;
    wire new_AGEMA_signal_98 ;
    wire new_AGEMA_signal_99 ;
    wire new_AGEMA_signal_100 ;
    wire new_AGEMA_signal_101 ;
    wire new_AGEMA_signal_102 ;
    wire new_AGEMA_signal_103 ;
    wire new_AGEMA_signal_104 ;
    wire new_AGEMA_signal_105 ;
    wire new_AGEMA_signal_106 ;
    wire new_AGEMA_signal_107 ;
    wire new_AGEMA_signal_108 ;
    wire new_AGEMA_signal_109 ;
    wire new_AGEMA_signal_110 ;
    wire new_AGEMA_signal_111 ;
    wire new_AGEMA_signal_112 ;
    wire new_AGEMA_signal_113 ;
    wire new_AGEMA_signal_114 ;
    wire new_AGEMA_signal_151 ;
    wire new_AGEMA_signal_152 ;
    wire new_AGEMA_signal_153 ;
    wire new_AGEMA_signal_154 ;
    wire new_AGEMA_signal_155 ;
    wire new_AGEMA_signal_156 ;
    wire new_AGEMA_signal_157 ;
    wire new_AGEMA_signal_158 ;
    wire new_AGEMA_signal_159 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_161 ;
    wire new_AGEMA_signal_162 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_166 ;
    wire new_AGEMA_signal_167 ;
    wire new_AGEMA_signal_168 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_171 ;
    wire new_AGEMA_signal_172 ;
    wire new_AGEMA_signal_173 ;
    wire new_AGEMA_signal_174 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_181 ;
    wire new_AGEMA_signal_182 ;
    wire new_AGEMA_signal_183 ;
    wire new_AGEMA_signal_184 ;
    wire new_AGEMA_signal_185 ;
    wire new_AGEMA_signal_186 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_191 ;
    wire new_AGEMA_signal_192 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) U5 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR_i1_U1 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .c ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, XX[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR_i2_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, XX[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR0_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, XX[2]}), .c ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, Q0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR1_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, XX[1]}), .c ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, Q1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) XOR3_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}), .c ({new_AGEMA_signal_66, new_AGEMA_signal_65, new_AGEMA_signal_64, Q4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR5_U1 ( .a ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, XX[2]}), .b ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}), .c ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, Q6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) XOR6_U1 ( .a ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, Q1}), .b ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, Q6}), .c ({new_AGEMA_signal_81, new_AGEMA_signal_80, new_AGEMA_signal_79, L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR8_U1 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}), .c ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, L2}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_26 ( .C (clk), .D (Q0), .Q (new_AGEMA_signal_151) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C (clk), .D (new_AGEMA_signal_58), .Q (new_AGEMA_signal_153) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C (clk), .D (new_AGEMA_signal_59), .Q (new_AGEMA_signal_155) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C (clk), .D (new_AGEMA_signal_60), .Q (new_AGEMA_signal_157) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C (clk), .D (L1), .Q (new_AGEMA_signal_159) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C (clk), .D (new_AGEMA_signal_79), .Q (new_AGEMA_signal_161) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C (clk), .D (new_AGEMA_signal_80), .Q (new_AGEMA_signal_163) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C (clk), .D (new_AGEMA_signal_81), .Q (new_AGEMA_signal_165) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C (clk), .D (XX[2]), .Q (new_AGEMA_signal_167) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C (clk), .D (new_AGEMA_signal_52), .Q (new_AGEMA_signal_169) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C (clk), .D (new_AGEMA_signal_53), .Q (new_AGEMA_signal_171) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C (clk), .D (new_AGEMA_signal_54), .Q (new_AGEMA_signal_173) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C (clk), .D (XX[1]), .Q (new_AGEMA_signal_175) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C (clk), .D (new_AGEMA_signal_46), .Q (new_AGEMA_signal_177) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C (clk), .D (new_AGEMA_signal_47), .Q (new_AGEMA_signal_179) ) ;
    buf_clk new_AGEMA_reg_buffer_56 ( .C (clk), .D (new_AGEMA_signal_48), .Q (new_AGEMA_signal_181) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C (clk), .D (X_s0[1]), .Q (new_AGEMA_signal_183) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C (clk), .D (X_s1[1]), .Q (new_AGEMA_signal_185) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C (clk), .D (X_s2[1]), .Q (new_AGEMA_signal_187) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C (clk), .D (X_s3[1]), .Q (new_AGEMA_signal_189) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C (clk), .D (Q6), .Q (new_AGEMA_signal_199) ) ;
    buf_clk new_AGEMA_reg_buffer_76 ( .C (clk), .D (new_AGEMA_signal_67), .Q (new_AGEMA_signal_201) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C (clk), .D (new_AGEMA_signal_68), .Q (new_AGEMA_signal_203) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C (clk), .D (new_AGEMA_signal_69), .Q (new_AGEMA_signal_205) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C (clk), .D (L2), .Q (new_AGEMA_signal_207) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C (clk), .D (new_AGEMA_signal_70), .Q (new_AGEMA_signal_211) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C (clk), .D (new_AGEMA_signal_71), .Q (new_AGEMA_signal_215) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C (clk), .D (new_AGEMA_signal_72), .Q (new_AGEMA_signal_219) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) AND1_U1 ( .a ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}), .b ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, Q1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, T0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR2_U1 ( .a ({new_AGEMA_signal_158, new_AGEMA_signal_156, new_AGEMA_signal_154, new_AGEMA_signal_152}), .b ({new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, T0}), .c ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, Q2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) AND3_U1 ( .a ({new_AGEMA_signal_42, new_AGEMA_signal_41, new_AGEMA_signal_40, n2}), .b ({new_AGEMA_signal_66, new_AGEMA_signal_65, new_AGEMA_signal_64, Q4}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR7_U1 ( .a ({new_AGEMA_signal_166, new_AGEMA_signal_164, new_AGEMA_signal_162, new_AGEMA_signal_160}), .b ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, T2}), .c ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, Q7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR11_U1 ( .a ({new_AGEMA_signal_174, new_AGEMA_signal_172, new_AGEMA_signal_170, new_AGEMA_signal_168}), .b ({new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, T0}), .c ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, L3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) XOR12_U1 ( .a ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, L3}), .b ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, T2}), .c ({new_AGEMA_signal_102, new_AGEMA_signal_101, new_AGEMA_signal_100, YY[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) XOR13_U1 ( .a ({new_AGEMA_signal_182, new_AGEMA_signal_180, new_AGEMA_signal_178, new_AGEMA_signal_176}), .b ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, T2}), .c ({new_AGEMA_signal_93, new_AGEMA_signal_92, new_AGEMA_signal_91, YY[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C (clk), .D (new_AGEMA_signal_151), .Q (new_AGEMA_signal_152) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C (clk), .D (new_AGEMA_signal_153), .Q (new_AGEMA_signal_154) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C (clk), .D (new_AGEMA_signal_155), .Q (new_AGEMA_signal_156) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C (clk), .D (new_AGEMA_signal_157), .Q (new_AGEMA_signal_158) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C (clk), .D (new_AGEMA_signal_159), .Q (new_AGEMA_signal_160) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C (clk), .D (new_AGEMA_signal_161), .Q (new_AGEMA_signal_162) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C (clk), .D (new_AGEMA_signal_163), .Q (new_AGEMA_signal_164) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C (clk), .D (new_AGEMA_signal_165), .Q (new_AGEMA_signal_166) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C (clk), .D (new_AGEMA_signal_167), .Q (new_AGEMA_signal_168) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C (clk), .D (new_AGEMA_signal_169), .Q (new_AGEMA_signal_170) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C (clk), .D (new_AGEMA_signal_171), .Q (new_AGEMA_signal_172) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C (clk), .D (new_AGEMA_signal_173), .Q (new_AGEMA_signal_174) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C (clk), .D (new_AGEMA_signal_175), .Q (new_AGEMA_signal_176) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C (clk), .D (new_AGEMA_signal_177), .Q (new_AGEMA_signal_178) ) ;
    buf_clk new_AGEMA_reg_buffer_55 ( .C (clk), .D (new_AGEMA_signal_179), .Q (new_AGEMA_signal_180) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C (clk), .D (new_AGEMA_signal_181), .Q (new_AGEMA_signal_182) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C (clk), .D (new_AGEMA_signal_183), .Q (new_AGEMA_signal_184) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C (clk), .D (new_AGEMA_signal_185), .Q (new_AGEMA_signal_186) ) ;
    buf_clk new_AGEMA_reg_buffer_63 ( .C (clk), .D (new_AGEMA_signal_187), .Q (new_AGEMA_signal_188) ) ;
    buf_clk new_AGEMA_reg_buffer_65 ( .C (clk), .D (new_AGEMA_signal_189), .Q (new_AGEMA_signal_190) ) ;
    buf_clk new_AGEMA_reg_buffer_75 ( .C (clk), .D (new_AGEMA_signal_199), .Q (new_AGEMA_signal_200) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C (clk), .D (new_AGEMA_signal_201), .Q (new_AGEMA_signal_202) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C (clk), .D (new_AGEMA_signal_203), .Q (new_AGEMA_signal_204) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C (clk), .D (new_AGEMA_signal_205), .Q (new_AGEMA_signal_206) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C (clk), .D (new_AGEMA_signal_207), .Q (new_AGEMA_signal_208) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C (clk), .D (new_AGEMA_signal_211), .Q (new_AGEMA_signal_212) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C (clk), .D (new_AGEMA_signal_215), .Q (new_AGEMA_signal_216) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C (clk), .D (new_AGEMA_signal_219), .Q (new_AGEMA_signal_220) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_66 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_191) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C (clk), .D (new_AGEMA_signal_76), .Q (new_AGEMA_signal_193) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C (clk), .D (new_AGEMA_signal_77), .Q (new_AGEMA_signal_195) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C (clk), .D (new_AGEMA_signal_78), .Q (new_AGEMA_signal_197) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C (clk), .D (new_AGEMA_signal_208), .Q (new_AGEMA_signal_209) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C (clk), .D (new_AGEMA_signal_212), .Q (new_AGEMA_signal_213) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C (clk), .D (new_AGEMA_signal_216), .Q (new_AGEMA_signal_217) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C (clk), .D (new_AGEMA_signal_220), .Q (new_AGEMA_signal_221) ) ;
    buf_clk new_AGEMA_reg_buffer_98 ( .C (clk), .D (L3), .Q (new_AGEMA_signal_223) ) ;
    buf_clk new_AGEMA_reg_buffer_100 ( .C (clk), .D (new_AGEMA_signal_88), .Q (new_AGEMA_signal_225) ) ;
    buf_clk new_AGEMA_reg_buffer_102 ( .C (clk), .D (new_AGEMA_signal_89), .Q (new_AGEMA_signal_227) ) ;
    buf_clk new_AGEMA_reg_buffer_104 ( .C (clk), .D (new_AGEMA_signal_90), .Q (new_AGEMA_signal_229) ) ;
    buf_clk new_AGEMA_reg_buffer_106 ( .C (clk), .D (YY[1]), .Q (new_AGEMA_signal_231) ) ;
    buf_clk new_AGEMA_reg_buffer_108 ( .C (clk), .D (new_AGEMA_signal_100), .Q (new_AGEMA_signal_233) ) ;
    buf_clk new_AGEMA_reg_buffer_110 ( .C (clk), .D (new_AGEMA_signal_101), .Q (new_AGEMA_signal_235) ) ;
    buf_clk new_AGEMA_reg_buffer_112 ( .C (clk), .D (new_AGEMA_signal_102), .Q (new_AGEMA_signal_237) ) ;
    buf_clk new_AGEMA_reg_buffer_114 ( .C (clk), .D (YY[0]), .Q (new_AGEMA_signal_239) ) ;
    buf_clk new_AGEMA_reg_buffer_116 ( .C (clk), .D (new_AGEMA_signal_91), .Q (new_AGEMA_signal_241) ) ;
    buf_clk new_AGEMA_reg_buffer_118 ( .C (clk), .D (new_AGEMA_signal_92), .Q (new_AGEMA_signal_243) ) ;
    buf_clk new_AGEMA_reg_buffer_120 ( .C (clk), .D (new_AGEMA_signal_93), .Q (new_AGEMA_signal_245) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) AND2_U1 ( .a ({new_AGEMA_signal_190, new_AGEMA_signal_188, new_AGEMA_signal_186, new_AGEMA_signal_184}), .b ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, Q2}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR4_U1 ( .a ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, T1}), .b ({new_AGEMA_signal_198, new_AGEMA_signal_196, new_AGEMA_signal_194, new_AGEMA_signal_192}), .c ({new_AGEMA_signal_105, new_AGEMA_signal_104, new_AGEMA_signal_103, L0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) AND4_U1 ( .a ({new_AGEMA_signal_206, new_AGEMA_signal_204, new_AGEMA_signal_202, new_AGEMA_signal_200}), .b ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, Q7}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR81_U1 ( .a ({new_AGEMA_signal_222, new_AGEMA_signal_218, new_AGEMA_signal_214, new_AGEMA_signal_210}), .b ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, T1}), .c ({new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, L2_T1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) XOR9_U1 ( .a ({new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, L2_T1}), .b ({new_AGEMA_signal_230, new_AGEMA_signal_228, new_AGEMA_signal_226, new_AGEMA_signal_224}), .c ({new_AGEMA_signal_111, new_AGEMA_signal_110, new_AGEMA_signal_109, YY[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) XOR10_U1 ( .a ({new_AGEMA_signal_105, new_AGEMA_signal_104, new_AGEMA_signal_103, L0}), .b ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, T3}), .c ({new_AGEMA_signal_114, new_AGEMA_signal_113, new_AGEMA_signal_112, YY[2]}) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C (clk), .D (new_AGEMA_signal_191), .Q (new_AGEMA_signal_192) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C (clk), .D (new_AGEMA_signal_193), .Q (new_AGEMA_signal_194) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C (clk), .D (new_AGEMA_signal_195), .Q (new_AGEMA_signal_196) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C (clk), .D (new_AGEMA_signal_197), .Q (new_AGEMA_signal_198) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C (clk), .D (new_AGEMA_signal_209), .Q (new_AGEMA_signal_210) ) ;
    buf_clk new_AGEMA_reg_buffer_89 ( .C (clk), .D (new_AGEMA_signal_213), .Q (new_AGEMA_signal_214) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C (clk), .D (new_AGEMA_signal_217), .Q (new_AGEMA_signal_218) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C (clk), .D (new_AGEMA_signal_221), .Q (new_AGEMA_signal_222) ) ;
    buf_clk new_AGEMA_reg_buffer_99 ( .C (clk), .D (new_AGEMA_signal_223), .Q (new_AGEMA_signal_224) ) ;
    buf_clk new_AGEMA_reg_buffer_101 ( .C (clk), .D (new_AGEMA_signal_225), .Q (new_AGEMA_signal_226) ) ;
    buf_clk new_AGEMA_reg_buffer_103 ( .C (clk), .D (new_AGEMA_signal_227), .Q (new_AGEMA_signal_228) ) ;
    buf_clk new_AGEMA_reg_buffer_105 ( .C (clk), .D (new_AGEMA_signal_229), .Q (new_AGEMA_signal_230) ) ;
    buf_clk new_AGEMA_reg_buffer_107 ( .C (clk), .D (new_AGEMA_signal_231), .Q (new_AGEMA_signal_232) ) ;
    buf_clk new_AGEMA_reg_buffer_109 ( .C (clk), .D (new_AGEMA_signal_233), .Q (new_AGEMA_signal_234) ) ;
    buf_clk new_AGEMA_reg_buffer_111 ( .C (clk), .D (new_AGEMA_signal_235), .Q (new_AGEMA_signal_236) ) ;
    buf_clk new_AGEMA_reg_buffer_113 ( .C (clk), .D (new_AGEMA_signal_237), .Q (new_AGEMA_signal_238) ) ;
    buf_clk new_AGEMA_reg_buffer_115 ( .C (clk), .D (new_AGEMA_signal_239), .Q (new_AGEMA_signal_240) ) ;
    buf_clk new_AGEMA_reg_buffer_117 ( .C (clk), .D (new_AGEMA_signal_241), .Q (new_AGEMA_signal_242) ) ;
    buf_clk new_AGEMA_reg_buffer_119 ( .C (clk), .D (new_AGEMA_signal_243), .Q (new_AGEMA_signal_244) ) ;
    buf_clk new_AGEMA_reg_buffer_121 ( .C (clk), .D (new_AGEMA_signal_245), .Q (new_AGEMA_signal_246) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_238, new_AGEMA_signal_236, new_AGEMA_signal_234, new_AGEMA_signal_232}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_246, new_AGEMA_signal_244, new_AGEMA_signal_242, new_AGEMA_signal_240}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_111, new_AGEMA_signal_110, new_AGEMA_signal_109, YY[3]}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_114, new_AGEMA_signal_113, new_AGEMA_signal_112, YY[2]}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
