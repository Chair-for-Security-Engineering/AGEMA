module Reg1(x, y);
 input [174:0] x;
 output [173:0] y;

  assign y[14] = x[3];
  assign y[15] = x[1];
  assign y[16] = x[2];
  assign y[17] = x[170];
  assign y[18] = x[99];
  assign y[19] = x[168];
  assign y[20] = x[169];
  assign y[21] = x[102];
  assign y[22] = x[103];
  assign y[23] = x[98];
  assign y[24] = x[100];
  assign y[25] = x[101];
  assign y[170] = x[171];
  assign y[171] = x[172];
  assign y[172] = x[173];
  assign y[173] = x[174];
  register_stage #(.WIDTH(158)) inst_0(.clk(x[0]), .D({x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[104],x[105],x[106],x[107],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[18],x[19],x[20],x[21],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169]}));
endmodule

module Reg2(x, y);
 input [315:0] x;
 output [314:0] y;

  assign y[70] = x[11];
  assign y[71] = x[12];
  assign y[72] = x[13];
  assign y[73] = x[14];
  assign y[74] = x[15];
  assign y[75] = x[1];
  assign y[76] = x[2];
  assign y[77] = x[3];
  assign y[78] = x[4];
  assign y[79] = x[5];
  assign y[80] = x[6];
  assign y[81] = x[7];
  assign y[82] = x[8];
  assign y[83] = x[9];
  assign y[84] = x[10];
  assign y[85] = x[306];
  assign y[86] = x[307];
  assign y[87] = x[308];
  assign y[88] = x[309];
  assign y[89] = x[310];
  assign y[90] = x[191];
  assign y[91] = x[192];
  assign y[92] = x[193];
  assign y[93] = x[194];
  assign y[94] = x[195];
  assign y[95] = x[296];
  assign y[96] = x[297];
  assign y[97] = x[298];
  assign y[98] = x[299];
  assign y[99] = x[300];
  assign y[100] = x[301];
  assign y[101] = x[302];
  assign y[102] = x[303];
  assign y[103] = x[304];
  assign y[104] = x[305];
  assign y[105] = x[206];
  assign y[106] = x[207];
  assign y[107] = x[208];
  assign y[108] = x[209];
  assign y[109] = x[210];
  assign y[110] = x[211];
  assign y[111] = x[212];
  assign y[112] = x[213];
  assign y[113] = x[214];
  assign y[114] = x[215];
  assign y[115] = x[186];
  assign y[116] = x[187];
  assign y[117] = x[188];
  assign y[118] = x[189];
  assign y[119] = x[190];
  assign y[120] = x[196];
  assign y[121] = x[197];
  assign y[122] = x[198];
  assign y[123] = x[199];
  assign y[124] = x[200];
  assign y[125] = x[201];
  assign y[126] = x[202];
  assign y[127] = x[203];
  assign y[128] = x[204];
  assign y[129] = x[205];
  assign y[310] = x[311];
  assign y[311] = x[312];
  assign y[312] = x[313];
  assign y[313] = x[314];
  assign y[314] = x[315];
  register_stage #(.WIDTH(250)) inst_0(.clk(x[0]), .D({x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[216],x[217],x[218],x[219],x[220],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[272],x[273],x[274],x[275],x[276],x[277],x[278],x[279],x[280],x[281],x[282],x[283],x[284],x[285],x[286],x[287],x[288],x[289],x[290],x[291],x[292],x[293],x[294],x[295],x[86],x[87],x[88],x[89],x[90],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272],y[273],y[274],y[275],y[276],y[277],y[278],y[279],y[280],y[281],y[282],y[283],y[284],y[285],y[286],y[287],y[288],y[289],y[290],y[291],y[292],y[293],y[294],y[295],y[296],y[297],y[298],y[299],y[300],y[301],y[302],y[303],y[304],y[305],y[306],y[307],y[308],y[309]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx266(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx267(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx268(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx269(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx270(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx271(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx272(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx273(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx274(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx275(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx276(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx277(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx278(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx279(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx280(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx281(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx282(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx283(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx284(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx285(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx286(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx287(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx288(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx289(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx290(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx291(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx292(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx293(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx294(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx295(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx296(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx297(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx298(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx299(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx300(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx301(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx302(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx303(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx304(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx305(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx306(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx307(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx308(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx309(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx310(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx311(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx312(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx313(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx314(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [410:0] x;
 output [236:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx29 Fx29_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx30 Fx30_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx34 Fx34_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx35 Fx35_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx39 Fx39_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx40 Fx40_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx44 Fx44_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx45 Fx45_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx49 Fx49_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx50 Fx50_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx54 Fx54_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx55 Fx55_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx59 Fx59_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx60 Fx60_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx64 Fx64_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx65 Fx65_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx69 Fx69_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx70 Fx70_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx74 Fx74_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx75 Fx75_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx79 Fx79_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx80 Fx80_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx84 Fx84_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx85 Fx85_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx89 Fx89_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx90 Fx90_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx94 Fx94_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx95 Fx95_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx99 Fx99_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx100 Fx100_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx104 Fx104_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx105 Fx105_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx109 Fx109_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx110 Fx110_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx114 Fx114_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx115 Fx115_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx119 Fx119_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx120 Fx120_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx124 Fx124_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx125 Fx125_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx129 Fx129_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx130 Fx130_inst(.x({x[82], x[81], x[80], x[79], x[78]}), .y(y[52]));
  Fx131 Fx131_inst(.x({x[83], x[81]}), .y(y[53]));
  Fx132 Fx132_inst(.x({x[84], x[80]}), .y(y[54]));
  Fx133 Fx133_inst(.x({x[85], x[79]}), .y(y[55]));
  Fx134 Fx134_inst(.x({x[86], x[78]}), .y(y[56]));
  Fx135 Fx135_inst(.x({x[91], x[90], x[89], x[88], x[87]}), .y(y[57]));
  Fx136 Fx136_inst(.x({x[92], x[90]}), .y(y[58]));
  Fx137 Fx137_inst(.x({x[93], x[89]}), .y(y[59]));
  Fx138 Fx138_inst(.x({x[94], x[88]}), .y(y[60]));
  Fx139 Fx139_inst(.x({x[95], x[87]}), .y(y[61]));
  Fx140 Fx140_inst(.x({x[100], x[99], x[98], x[97], x[96]}), .y(y[62]));
  Fx141 Fx141_inst(.x({x[101], x[99]}), .y(y[63]));
  Fx142 Fx142_inst(.x({x[102], x[98]}), .y(y[64]));
  Fx143 Fx143_inst(.x({x[103], x[97]}), .y(y[65]));
  Fx144 Fx144_inst(.x({x[104], x[96]}), .y(y[66]));
  Fx145 Fx145_inst(.x({x[109], x[108], x[107], x[106], x[105]}), .y(y[67]));
  Fx146 Fx146_inst(.x({x[110], x[108]}), .y(y[68]));
  Fx147 Fx147_inst(.x({x[111], x[107]}), .y(y[69]));
  Fx148 Fx148_inst(.x({x[112], x[106]}), .y(y[70]));
  Fx149 Fx149_inst(.x({x[113], x[105]}), .y(y[71]));
  Fx150 Fx150_inst(.x({x[118], x[117], x[116], x[115], x[114]}), .y(y[72]));
  Fx151 Fx151_inst(.x({x[119], x[117]}), .y(y[73]));
  Fx152 Fx152_inst(.x({x[120], x[116]}), .y(y[74]));
  Fx153 Fx153_inst(.x({x[121], x[115]}), .y(y[75]));
  Fx154 Fx154_inst(.x({x[122], x[114]}), .y(y[76]));
  Fx155 Fx155_inst(.x({x[127], x[126], x[125], x[124], x[123]}), .y(y[77]));
  Fx156 Fx156_inst(.x({x[128], x[126]}), .y(y[78]));
  Fx157 Fx157_inst(.x({x[129], x[125]}), .y(y[79]));
  Fx158 Fx158_inst(.x({x[130], x[124]}), .y(y[80]));
  Fx159 Fx159_inst(.x({x[131], x[123]}), .y(y[81]));
  Fx160 Fx160_inst(.x({x[136], x[135], x[134], x[133], x[132]}), .y(y[82]));
  Fx161 Fx161_inst(.x({x[137], x[135]}), .y(y[83]));
  Fx162 Fx162_inst(.x({x[138], x[134]}), .y(y[84]));
  Fx163 Fx163_inst(.x({x[139], x[133]}), .y(y[85]));
  Fx164 Fx164_inst(.x({x[140], x[132]}), .y(y[86]));
  Fx165 Fx165_inst(.x({x[145], x[144], x[143], x[142], x[141]}), .y(y[87]));
  Fx166 Fx166_inst(.x({x[146], x[144]}), .y(y[88]));
  Fx167 Fx167_inst(.x({x[147], x[143]}), .y(y[89]));
  Fx168 Fx168_inst(.x({x[148], x[142]}), .y(y[90]));
  Fx169 Fx169_inst(.x({x[149], x[141]}), .y(y[91]));
  Fx170 Fx170_inst(.x({x[154], x[153], x[152], x[151], x[150]}), .y(y[92]));
  Fx171 Fx171_inst(.x({x[155], x[153]}), .y(y[93]));
  Fx172 Fx172_inst(.x({x[156], x[152]}), .y(y[94]));
  Fx173 Fx173_inst(.x({x[157], x[151]}), .y(y[95]));
  Fx174 Fx174_inst(.x({x[158], x[150]}), .y(y[96]));
  Fx175 Fx175_inst(.x({x[163], x[162], x[161], x[160], x[159]}), .y(y[97]));
  Fx176 Fx176_inst(.x({x[164], x[162]}), .y(y[98]));
  Fx177 Fx177_inst(.x({x[165], x[161]}), .y(y[99]));
  Fx178 Fx178_inst(.x({x[166], x[160]}), .y(y[100]));
  Fx179 Fx179_inst(.x({x[167], x[159]}), .y(y[101]));
  Fx180 Fx180_inst(.x({x[172], x[171], x[170], x[169], x[168]}), .y(y[102]));
  Fx181 Fx181_inst(.x({x[173], x[171]}), .y(y[103]));
  Fx182 Fx182_inst(.x({x[174], x[170]}), .y(y[104]));
  Fx183 Fx183_inst(.x({x[175], x[169]}), .y(y[105]));
  Fx184 Fx184_inst(.x({x[176], x[168]}), .y(y[106]));
  Fx185 Fx185_inst(.x({x[181], x[180], x[179], x[178], x[177]}), .y(y[107]));
  Fx186 Fx186_inst(.x({x[182], x[180]}), .y(y[108]));
  Fx187 Fx187_inst(.x({x[183], x[179]}), .y(y[109]));
  Fx188 Fx188_inst(.x({x[184], x[178]}), .y(y[110]));
  Fx189 Fx189_inst(.x({x[185], x[177]}), .y(y[111]));
  Fx190 Fx190_inst(.x({x[190], x[189], x[188], x[187], x[186]}), .y(y[112]));
  Fx191 Fx191_inst(.x({x[191], x[189]}), .y(y[113]));
  Fx192 Fx192_inst(.x({x[192], x[188]}), .y(y[114]));
  Fx193 Fx193_inst(.x({x[193], x[187]}), .y(y[115]));
  Fx194 Fx194_inst(.x({x[194], x[186]}), .y(y[116]));
  Fx195 Fx195_inst(.x({x[199], x[198], x[197], x[196], x[195]}), .y(y[117]));
  Fx196 Fx196_inst(.x({x[200], x[198]}), .y(y[118]));
  Fx197 Fx197_inst(.x({x[201], x[197]}), .y(y[119]));
  Fx198 Fx198_inst(.x({x[202], x[196]}), .y(y[120]));
  Fx199 Fx199_inst(.x({x[203], x[195]}), .y(y[121]));
  Fx200 Fx200_inst(.x({x[208], x[207], x[206], x[205], x[204]}), .y(y[122]));
  Fx201 Fx201_inst(.x({x[209], x[207]}), .y(y[123]));
  Fx202 Fx202_inst(.x({x[210], x[206]}), .y(y[124]));
  Fx203 Fx203_inst(.x({x[211], x[205]}), .y(y[125]));
  Fx204 Fx204_inst(.x({x[212], x[204]}), .y(y[126]));
  Fx205 Fx205_inst(.x({x[217], x[216], x[215], x[214], x[213]}), .y(y[127]));
  Fx206 Fx206_inst(.x({x[218], x[216]}), .y(y[128]));
  Fx207 Fx207_inst(.x({x[219], x[215]}), .y(y[129]));
  Fx208 Fx208_inst(.x({x[220], x[214]}), .y(y[130]));
  Fx209 Fx209_inst(.x({x[221], x[213]}), .y(y[131]));
  Fx210 Fx210_inst(.x({x[226], x[225], x[224], x[223], x[222]}), .y(y[132]));
  Fx211 Fx211_inst(.x({x[227], x[225]}), .y(y[133]));
  Fx212 Fx212_inst(.x({x[228], x[224]}), .y(y[134]));
  Fx213 Fx213_inst(.x({x[229], x[223]}), .y(y[135]));
  Fx214 Fx214_inst(.x({x[230], x[222]}), .y(y[136]));
  Fx215 Fx215_inst(.x({x[235], x[234], x[233], x[232], x[231]}), .y(y[137]));
  Fx216 Fx216_inst(.x({x[236], x[234]}), .y(y[138]));
  Fx217 Fx217_inst(.x({x[237], x[233]}), .y(y[139]));
  Fx218 Fx218_inst(.x({x[238], x[232]}), .y(y[140]));
  Fx219 Fx219_inst(.x({x[239], x[231]}), .y(y[141]));
  Fx220 Fx220_inst(.x({x[244], x[243], x[242], x[241], x[240]}), .y(y[142]));
  Fx221 Fx221_inst(.x({x[245], x[243]}), .y(y[143]));
  Fx222 Fx222_inst(.x({x[246], x[242]}), .y(y[144]));
  Fx223 Fx223_inst(.x({x[247], x[241]}), .y(y[145]));
  Fx224 Fx224_inst(.x({x[248], x[240]}), .y(y[146]));
  Fx225 Fx225_inst(.x({x[253], x[252], x[251], x[250], x[249]}), .y(y[147]));
  Fx226 Fx226_inst(.x({x[254], x[252]}), .y(y[148]));
  Fx227 Fx227_inst(.x({x[255], x[251]}), .y(y[149]));
  Fx228 Fx228_inst(.x({x[256], x[250]}), .y(y[150]));
  Fx229 Fx229_inst(.x({x[257], x[249]}), .y(y[151]));
  Fx230 Fx230_inst(.x({x[262], x[261], x[260], x[259], x[258]}), .y(y[152]));
  Fx231 Fx231_inst(.x({x[263], x[261]}), .y(y[153]));
  Fx232 Fx232_inst(.x({x[264], x[260]}), .y(y[154]));
  Fx233 Fx233_inst(.x({x[265], x[259]}), .y(y[155]));
  Fx234 Fx234_inst(.x({x[266], x[258]}), .y(y[156]));
  Fx235 Fx235_inst(.x({x[271], x[270], x[269], x[268], x[267]}), .y(y[157]));
  Fx236 Fx236_inst(.x({x[272], x[270]}), .y(y[158]));
  Fx237 Fx237_inst(.x({x[273], x[269]}), .y(y[159]));
  Fx238 Fx238_inst(.x({x[274], x[268]}), .y(y[160]));
  Fx239 Fx239_inst(.x({x[275], x[267]}), .y(y[161]));
  Fx240 Fx240_inst(.x({x[280], x[279], x[278], x[277], x[276]}), .y(y[162]));
  Fx241 Fx241_inst(.x({x[281], x[279]}), .y(y[163]));
  Fx242 Fx242_inst(.x({x[282], x[278]}), .y(y[164]));
  Fx243 Fx243_inst(.x({x[283], x[277]}), .y(y[165]));
  Fx244 Fx244_inst(.x({x[284], x[276]}), .y(y[166]));
  Fx245 Fx245_inst(.x({x[289], x[288], x[287], x[286], x[285]}), .y(y[167]));
  Fx246 Fx246_inst(.x({x[290], x[288]}), .y(y[168]));
  Fx247 Fx247_inst(.x({x[291], x[287]}), .y(y[169]));
  Fx248 Fx248_inst(.x({x[292], x[286]}), .y(y[170]));
  Fx249 Fx249_inst(.x({x[293], x[285]}), .y(y[171]));
  Fx250 Fx250_inst(.x({x[298], x[297], x[296], x[295], x[294]}), .y(y[172]));
  Fx251 Fx251_inst(.x({x[299], x[297]}), .y(y[173]));
  Fx252 Fx252_inst(.x({x[300], x[296]}), .y(y[174]));
  Fx253 Fx253_inst(.x({x[301], x[295]}), .y(y[175]));
  Fx254 Fx254_inst(.x({x[302], x[294]}), .y(y[176]));
  Fx255 Fx255_inst(.x({x[307], x[306], x[305], x[304], x[303]}), .y(y[177]));
  Fx256 Fx256_inst(.x({x[308], x[306]}), .y(y[178]));
  Fx257 Fx257_inst(.x({x[309], x[305]}), .y(y[179]));
  Fx258 Fx258_inst(.x({x[310], x[304]}), .y(y[180]));
  Fx259 Fx259_inst(.x({x[311], x[303]}), .y(y[181]));
  Fx260 Fx260_inst(.x({x[316], x[315], x[314], x[313], x[312]}), .y(y[182]));
  Fx261 Fx261_inst(.x({x[317], x[315]}), .y(y[183]));
  Fx262 Fx262_inst(.x({x[318], x[314]}), .y(y[184]));
  Fx263 Fx263_inst(.x({x[319], x[313]}), .y(y[185]));
  Fx264 Fx264_inst(.x({x[320], x[312]}), .y(y[186]));
  Fx265 Fx265_inst(.x({x[325], x[324], x[323], x[322], x[321]}), .y(y[187]));
  Fx266 Fx266_inst(.x({x[326], x[324]}), .y(y[188]));
  Fx267 Fx267_inst(.x({x[327], x[323]}), .y(y[189]));
  Fx268 Fx268_inst(.x({x[328], x[322]}), .y(y[190]));
  Fx269 Fx269_inst(.x({x[329], x[321]}), .y(y[191]));
  Fx270 Fx270_inst(.x({x[334], x[333], x[332], x[331], x[330]}), .y(y[192]));
  Fx271 Fx271_inst(.x({x[335], x[333]}), .y(y[193]));
  Fx272 Fx272_inst(.x({x[336], x[332]}), .y(y[194]));
  Fx273 Fx273_inst(.x({x[337], x[331]}), .y(y[195]));
  Fx274 Fx274_inst(.x({x[338], x[330]}), .y(y[196]));
  Fx275 Fx275_inst(.x({x[343], x[342], x[341], x[340], x[339]}), .y(y[197]));
  Fx276 Fx276_inst(.x({x[344], x[342]}), .y(y[198]));
  Fx277 Fx277_inst(.x({x[345], x[341]}), .y(y[199]));
  Fx278 Fx278_inst(.x({x[346], x[340]}), .y(y[200]));
  Fx279 Fx279_inst(.x({x[347], x[339]}), .y(y[201]));
  Fx280 Fx280_inst(.x({x[352], x[351], x[350], x[349], x[348]}), .y(y[202]));
  Fx281 Fx281_inst(.x({x[353], x[351]}), .y(y[203]));
  Fx282 Fx282_inst(.x({x[354], x[350]}), .y(y[204]));
  Fx283 Fx283_inst(.x({x[355], x[349]}), .y(y[205]));
  Fx284 Fx284_inst(.x({x[356], x[348]}), .y(y[206]));
  Fx285 Fx285_inst(.x({x[361], x[360], x[359], x[358], x[357]}), .y(y[207]));
  Fx286 Fx286_inst(.x({x[362], x[360]}), .y(y[208]));
  Fx287 Fx287_inst(.x({x[363], x[359]}), .y(y[209]));
  Fx288 Fx288_inst(.x({x[364], x[358]}), .y(y[210]));
  Fx289 Fx289_inst(.x({x[365], x[357]}), .y(y[211]));
  Fx290 Fx290_inst(.x({x[370], x[369], x[368], x[367], x[366]}), .y(y[212]));
  Fx291 Fx291_inst(.x({x[371], x[369]}), .y(y[213]));
  Fx292 Fx292_inst(.x({x[372], x[368]}), .y(y[214]));
  Fx293 Fx293_inst(.x({x[373], x[367]}), .y(y[215]));
  Fx294 Fx294_inst(.x({x[374], x[366]}), .y(y[216]));
  Fx295 Fx295_inst(.x({x[379], x[378], x[377], x[376], x[375]}), .y(y[217]));
  Fx296 Fx296_inst(.x({x[380], x[378]}), .y(y[218]));
  Fx297 Fx297_inst(.x({x[381], x[377]}), .y(y[219]));
  Fx298 Fx298_inst(.x({x[382], x[376]}), .y(y[220]));
  Fx299 Fx299_inst(.x({x[383], x[375]}), .y(y[221]));
  Fx300 Fx300_inst(.x({x[388], x[387], x[386], x[385], x[384]}), .y(y[222]));
  Fx301 Fx301_inst(.x({x[389], x[387]}), .y(y[223]));
  Fx302 Fx302_inst(.x({x[390], x[386]}), .y(y[224]));
  Fx303 Fx303_inst(.x({x[391], x[385]}), .y(y[225]));
  Fx304 Fx304_inst(.x({x[392], x[384]}), .y(y[226]));
  Fx305 Fx305_inst(.x({x[397], x[396], x[395], x[394], x[393]}), .y(y[227]));
  Fx306 Fx306_inst(.x({x[398], x[396]}), .y(y[228]));
  Fx307 Fx307_inst(.x({x[399], x[395]}), .y(y[229]));
  Fx308 Fx308_inst(.x({x[400], x[394]}), .y(y[230]));
  Fx309 Fx309_inst(.x({x[401], x[393]}), .y(y[231]));
  Fx310 Fx310_inst(.x({x[406], x[405], x[404], x[403], x[402]}), .y(y[232]));
  Fx311 Fx311_inst(.x({x[407], x[405]}), .y(y[233]));
  Fx312 Fx312_inst(.x({x[408], x[404]}), .y(y[234]));
  Fx313 Fx313_inst(.x({x[409], x[403]}), .y(y[235]));
  Fx314 Fx314_inst(.x({x[410], x[402]}), .y(y[236]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [26:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[19] ^ x[8];
  assign t[11] = t[20] ^ x[11];
  assign t[12] = t[21] ^ x[14];
  assign t[13] = t[22] ^ x[17];
  assign t[14] = t[23] ^ x[20];
  assign t[15] = t[24] ^ x[23];
  assign t[16] = t[25] ^ x[26];
  assign t[17] = (x[0] & x[1]);
  assign t[18] = (x[3] & x[4]);
  assign t[19] = (x[6] & x[7]);
  assign t[1] = ~(t[8] & t[4]);
  assign t[20] = (x[9] & x[10]);
  assign t[21] = (x[12] & x[13]);
  assign t[22] = (x[15] & x[16]);
  assign t[23] = (x[18] & x[19]);
  assign t[24] = (x[21] & x[22]);
  assign t[25] = (x[24] & x[25]);
  assign t[2] = ~(t[9] | t[10]);
  assign t[3] = ~(t[5] | t[11]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13] & t[14]);
  assign t[7] = ~(t[15] & t[16]);
  assign t[8] = t[17] ^ x[2];
  assign t[9] = t[18] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind66(x, y);
 input [22:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[17] ^ t[18]);
  assign t[11] = ~(t[19]);
  assign t[12] = t[20] ^ x[2];
  assign t[13] = t[21] ^ x[5];
  assign t[14] = t[22] ^ x[8];
  assign t[15] = t[23] ^ x[11];
  assign t[16] = t[24] ^ x[16];
  assign t[17] = t[25] ^ x[18];
  assign t[18] = t[26] ^ x[20];
  assign t[19] = t[27] ^ x[22];
  assign t[1] = ~(t[5] & t[12]);
  assign t[20] = (x[0] & x[1]);
  assign t[21] = (x[3] & x[4]);
  assign t[22] = (x[6] & x[7]);
  assign t[23] = (x[9] & x[10]);
  assign t[24] = (x[14] & x[15]);
  assign t[25] = (x[14] & x[17]);
  assign t[26] = (x[14] & x[19]);
  assign t[27] = (x[14] & x[21]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[13]);
  assign t[4] = ~(t[14] & t[7]);
  assign t[5] = ~(t[14] | t[6]);
  assign t[6] = ~(t[15]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] ^ t[10]);
  assign t[9] = ~(t[11] | t[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind67(x, y);
 input [22:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[13]);
  assign t[12] = t[23] ? t[16] : t[24];
  assign t[13] = ~(t[25]);
  assign t[14] = ~(t[23] ^ t[26]);
  assign t[15] = ~(t[23] | t[26]);
  assign t[16] = ~(t[24] & t[17]);
  assign t[17] = ~(t[18] & t[13]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[5] & t[19]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = t[31] ^ x[16];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[20];
  assign t[26] = t[34] ^ x[22];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[14] & x[17]);
  assign t[33] = (x[14] & x[19]);
  assign t[34] = (x[14] & x[21]);
  assign t[3] = ~(t[20]);
  assign t[4] = ~(t[21] & t[7]);
  assign t[5] = ~(t[21] | t[6]);
  assign t[6] = ~(t[22]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] | t[10]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind68(x, y);
 input [22:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[27] | t[15]);
  assign t[12] = ~(t[28] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = t[29] ? t[12] : t[28];
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[18]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[27]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~(t[5] & t[23]);
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[28]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[16];
  assign t[28] = t[36] ^ x[18];
  assign t[29] = t[37] ^ x[20];
  assign t[2] = ~(t[6]);
  assign t[30] = t[38] ^ x[22];
  assign t[31] = (x[0] & x[1]);
  assign t[32] = (x[3] & x[4]);
  assign t[33] = (x[6] & x[7]);
  assign t[34] = (x[9] & x[10]);
  assign t[35] = (x[14] & x[15]);
  assign t[36] = (x[14] & x[17]);
  assign t[37] = (x[14] & x[19]);
  assign t[38] = (x[14] & x[21]);
  assign t[3] = ~(t[24]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[5] = ~(t[25] | t[6]);
  assign t[6] = ~(t[26]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind69(x, y);
 input [22:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[24] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[23] | t[25]);
  assign t[14] = ~(t[24]);
  assign t[15] = ~(t[18] & t[16]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[18] & t[14]);
  assign t[18] = ~(t[25]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[5] & t[19]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = t[31] ^ x[16];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[20];
  assign t[26] = t[34] ^ x[22];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[14] & x[17]);
  assign t[33] = (x[14] & x[19]);
  assign t[34] = (x[14] & x[21]);
  assign t[3] = ~(t[20]);
  assign t[4] = ~(t[21] & t[7]);
  assign t[5] = ~(t[21] | t[6]);
  assign t[6] = ~(t[22]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = t[23] ? t[12] : t[11];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind70(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind71(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind72(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind73(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind74(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind75(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind76(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind77(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind78(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind79(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind80(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind81(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind82(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind83(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind84(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind85(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind86(x, y);
 input [15:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[14];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[6] & x[13]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[15] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind87(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind88(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind89(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind90(x, y);
 input [15:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[14];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[6] & x[13]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[15] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind91(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind92(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind93(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind94(x, y);
 input [15:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[14];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[6] & x[13]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[15] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind95(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind96(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind97(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind98(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind99(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind100(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind101(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind102(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind103(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind104(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind105(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind106(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind107(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind108(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind109(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind110(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind111(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind112(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind113(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind114(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind115(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind116(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind117(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind118(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind119(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind120(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind121(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind122(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind123(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind124(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind125(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind126(x, y);
 input [18:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[18];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[3] & x[17]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind127(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind128(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind129(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind130(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind131(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind132(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind133(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind134(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[3] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind135(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind136(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind137(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind138(x, y);
 input [15:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[14];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[6] & x[13]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[15] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind139(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind140(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind141(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind142(x, y);
 input [15:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[14];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[6] & x[13]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[15] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind143(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind144(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind145(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind146(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind147(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind148(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[14];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[0] & x[13]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[15] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind149(x, y);
 input [13:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[12] : t[11];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind150(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind151(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind152(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind153(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind154(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind155(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind156(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind157(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind158(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind159(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind160(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind161(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind162(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind163(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind164(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind165(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind166(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind167(x, y);
 input [15:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[13];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[3] & x[12]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[14] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[15]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind168(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[12] : t[11];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[13]);
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind169(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind170(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind171(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind172(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind173(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind174(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind175(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind176(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind177(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind178(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind179(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind180(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind181(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind182(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind183(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind184(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind185(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind186(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[13];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[0] & x[12]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[14] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[15]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind187(x, y);
 input [13:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[12] : t[11];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind188(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind189(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind190(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind191(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind192(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind193(x, y);
 input [15:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[13];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[3] & x[12]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[14] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[15]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind194(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind195(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind196(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind197(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind198(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind199(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind200(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind201(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind202(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind203(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind204(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind205(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind206(x, y);
 input [28:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[15] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[21]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[13] = ~(x[26]);
  assign t[14] = ~(t[24]);
  assign t[15] = t[25] ^ x[2];
  assign t[16] = t[26] ^ x[5];
  assign t[17] = t[27] ^ x[8];
  assign t[18] = t[28] ^ x[11];
  assign t[19] = t[29] ^ x[15];
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = t[30] ^ x[18];
  assign t[21] = t[31] ^ x[21];
  assign t[22] = t[32] ^ x[23];
  assign t[23] = t[33] ^ x[25];
  assign t[24] = t[34] ^ x[28];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[16]);
  assign t[30] = (x[16] & x[17]);
  assign t[31] = (x[19] & x[20]);
  assign t[32] = (x[19] & x[22]);
  assign t[33] = (x[19] & x[24]);
  assign t[34] = (x[19] & x[27]);
  assign t[3] = ~(t[17] & t[6]);
  assign t[4] = ~(t[17] | t[7]);
  assign t[5] = t[18] ? t[9] : t[8];
  assign t[6] = t[10] ? x[12] : t[16];
  assign t[7] = ~(t[15]);
  assign t[8] = ~(t[11] ^ t[12]);
  assign t[9] = t[19] ^ t[20];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind207(x, y);
 input [31:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[22] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(x[22]);
  assign t[14] = ~(t[18] | t[16]);
  assign t[15] = t[29] ? t[19] : t[30];
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[29] ^ t[32]);
  assign t[18] = ~(t[29] | t[32]);
  assign t[19] = ~(t[30] & t[20]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[21] & t[16]);
  assign t[21] = ~(t[32]);
  assign t[22] = t[33] ^ x[2];
  assign t[23] = t[34] ^ x[5];
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[11];
  assign t[26] = t[37] ^ x[14];
  assign t[27] = t[38] ^ x[18];
  assign t[28] = t[39] ^ x[21];
  assign t[29] = t[40] ^ x[25];
  assign t[2] = ~(t[23]);
  assign t[30] = t[41] ^ x[27];
  assign t[31] = t[42] ^ x[29];
  assign t[32] = t[43] ^ x[31];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[6] & x[7]);
  assign t[36] = (x[9] & x[10]);
  assign t[37] = (x[12] & x[13]);
  assign t[38] = (x[16] & x[17]);
  assign t[39] = (x[19] & x[20]);
  assign t[3] = ~(t[24] & t[6]);
  assign t[40] = (x[23] & x[24]);
  assign t[41] = (x[23] & x[26]);
  assign t[42] = (x[23] & x[28]);
  assign t[43] = (x[23] & x[30]);
  assign t[4] = ~(t[24] | t[7]);
  assign t[5] = t[25] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[26];
  assign t[7] = ~(t[22]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = t[27] ^ t[28];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind208(x, y);
 input [31:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[26] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(x[22]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[34] & t[19]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = t[35] ? t[15] : t[34];
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[21]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[35] | t[36]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[34]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[8];
  assign t[29] = t[40] ^ x[11];
  assign t[2] = ~(t[27]);
  assign t[30] = t[41] ^ x[14];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[25];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[29];
  assign t[36] = t[47] ^ x[31];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[28] & t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[12] & x[13]);
  assign t[42] = (x[16] & x[17]);
  assign t[43] = (x[19] & x[20]);
  assign t[44] = (x[23] & x[24]);
  assign t[45] = (x[23] & x[26]);
  assign t[46] = (x[23] & x[28]);
  assign t[47] = (x[23] & x[30]);
  assign t[4] = ~(t[28] | t[7]);
  assign t[5] = t[29] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[30];
  assign t[7] = ~(t[26]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[31] ^ t[32];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind209(x, y);
 input [31:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[22] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = t[29] ? t[15] : t[14];
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(x[25]);
  assign t[14] = ~(t[30] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[29] | t[31]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[21] & t[19]);
  assign t[19] = ~(t[32]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[21] & t[17]);
  assign t[21] = ~(t[31]);
  assign t[22] = t[33] ^ x[2];
  assign t[23] = t[34] ^ x[5];
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[11];
  assign t[26] = t[37] ^ x[14];
  assign t[27] = t[38] ^ x[18];
  assign t[28] = t[39] ^ x[21];
  assign t[29] = t[40] ^ x[24];
  assign t[2] = ~(t[23]);
  assign t[30] = t[41] ^ x[27];
  assign t[31] = t[42] ^ x[29];
  assign t[32] = t[43] ^ x[31];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[6] & x[7]);
  assign t[36] = (x[9] & x[10]);
  assign t[37] = (x[12] & x[13]);
  assign t[38] = (x[16] & x[17]);
  assign t[39] = (x[19] & x[20]);
  assign t[3] = ~(t[24] & t[6]);
  assign t[40] = (x[22] & x[23]);
  assign t[41] = (x[22] & x[26]);
  assign t[42] = (x[22] & x[28]);
  assign t[43] = (x[22] & x[30]);
  assign t[4] = ~(t[24] | t[7]);
  assign t[5] = t[25] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[26];
  assign t[7] = ~(t[22]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[27] ^ t[28];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind210(x, y);
 input [24:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[18] ^ x[3];
  assign t[11] = t[19] ^ x[6];
  assign t[12] = t[20] ^ x[9];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[15];
  assign t[15] = t[23] ^ x[18];
  assign t[16] = t[24] ^ x[21];
  assign t[17] = t[25] ^ x[24];
  assign t[18] = (x[1] & x[2]);
  assign t[19] = (x[4] & x[5]);
  assign t[1] = ~(x[0]);
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[24] = (x[19] & x[20]);
  assign t[25] = (x[22] & x[23]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[7] & t[11];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14] & t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = t[0] & t[1];
endmodule

module R1ind211(x, y);
 input [29:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[16] ^ t[2]);
  assign t[10] = ~(t[21] | t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[22]);
  assign t[14] = t[15] & t[23];
  assign t[15] = ~(t[24] | t[25]);
  assign t[16] = t[26] ^ x[2];
  assign t[17] = t[27] ^ x[5];
  assign t[18] = t[28] ^ x[8];
  assign t[19] = t[29] ^ x[11];
  assign t[1] = ~(t[3]);
  assign t[20] = t[30] ^ x[14];
  assign t[21] = t[31] ^ x[17];
  assign t[22] = t[32] ^ x[20];
  assign t[23] = t[33] ^ x[23];
  assign t[24] = t[34] ^ x[26];
  assign t[25] = t[35] ^ x[29];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[3] & x[4]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[9] & x[10]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = (x[12] & x[13]);
  assign t[31] = (x[15] & x[16]);
  assign t[32] = (x[18] & x[19]);
  assign t[33] = (x[21] & x[22]);
  assign t[34] = (x[24] & x[25]);
  assign t[35] = (x[27] & x[28]);
  assign t[3] = ~(t[17]);
  assign t[4] = ~(t[18]);
  assign t[5] = ~(t[6] & t[19]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[20]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind212(x, y);
 input [26:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[19]);
  assign t[12] = t[13] & t[20];
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = t[23] ^ x[2];
  assign t[15] = t[24] ^ x[5];
  assign t[16] = t[25] ^ x[8];
  assign t[17] = t[26] ^ x[11];
  assign t[18] = t[27] ^ x[14];
  assign t[19] = t[28] ^ x[17];
  assign t[1] = t[14] ^ t[3];
  assign t[20] = t[29] ^ x[20];
  assign t[21] = t[30] ^ x[23];
  assign t[22] = t[31] ^ x[26];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[15] & x[16]);
  assign t[29] = (x[18] & x[19]);
  assign t[2] = ~(t[15]);
  assign t[30] = (x[21] & x[22]);
  assign t[31] = (x[24] & x[25]);
  assign t[3] = ~(t[4] & t[16]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[17]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[18] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind213(x, y);
 input [23:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] ^ t[13]);
  assign t[10] = ~(t[17]);
  assign t[11] = t[12] & t[18];
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[5];
  assign t[15] = t[23] ^ x[8];
  assign t[16] = t[24] ^ x[11];
  assign t[17] = t[25] ^ x[14];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[20];
  assign t[1] = ~(t[3]);
  assign t[20] = t[28] ^ x[23];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[3] & x[4]);
  assign t[23] = (x[6] & x[7]);
  assign t[24] = (x[9] & x[10]);
  assign t[25] = (x[12] & x[13]);
  assign t[26] = (x[15] & x[16]);
  assign t[27] = (x[18] & x[19]);
  assign t[28] = (x[21] & x[22]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[14]);
  assign t[4] = ~(t[15]);
  assign t[5] = ~(t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[16] | t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind214(x, y);
 input [20:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = t[18] ^ x[2];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[8];
  assign t[14] = t[21] ^ x[11];
  assign t[15] = t[22] ^ x[14];
  assign t[16] = t[23] ^ x[17];
  assign t[17] = t[24] ^ x[20];
  assign t[18] = (x[0] & x[1]);
  assign t[19] = (x[3] & x[4]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (x[6] & x[7]);
  assign t[21] = (x[9] & x[10]);
  assign t[22] = (x[12] & x[13]);
  assign t[23] = (x[15] & x[16]);
  assign t[24] = (x[18] & x[19]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[5]);
  assign t[5] = ~(t[13] | t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[10] & t[15];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind215(x, y);
 input [39:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[11] & t[24]);
  assign t[11] = t[25] & t[12];
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17]);
  assign t[15] = ~(t[26]);
  assign t[16] = t[18] & t[27];
  assign t[17] = ~(t[19] | t[20]);
  assign t[18] = ~(t[28] | t[29]);
  assign t[19] = ~(t[30] & t[31]);
  assign t[1] = t[21] ? t[4] : t[3];
  assign t[20] = ~(t[32] & t[33]);
  assign t[21] = t[34] ^ x[2];
  assign t[22] = t[35] ^ x[6];
  assign t[23] = t[36] ^ x[9];
  assign t[24] = t[37] ^ x[12];
  assign t[25] = t[38] ^ x[15];
  assign t[26] = t[39] ^ x[18];
  assign t[27] = t[40] ^ x[21];
  assign t[28] = t[41] ^ x[24];
  assign t[29] = t[42] ^ x[27];
  assign t[2] = ~(x[3]);
  assign t[30] = t[43] ^ x[30];
  assign t[31] = t[44] ^ x[33];
  assign t[32] = t[45] ^ x[36];
  assign t[33] = t[46] ^ x[39];
  assign t[34] = (x[0] & x[1]);
  assign t[35] = (x[4] & x[5]);
  assign t[36] = (x[7] & x[8]);
  assign t[37] = (x[10] & x[11]);
  assign t[38] = (x[13] & x[14]);
  assign t[39] = (x[16] & x[17]);
  assign t[3] = t[5] | t[6];
  assign t[40] = (x[19] & x[20]);
  assign t[41] = (x[22] & x[23]);
  assign t[42] = (x[25] & x[26]);
  assign t[43] = (x[28] & x[29]);
  assign t[44] = (x[31] & x[32]);
  assign t[45] = (x[34] & x[35]);
  assign t[46] = (x[37] & x[38]);
  assign t[4] = ~(t[5] | t[7]);
  assign t[5] = ~(t[22]);
  assign t[6] = ~(t[8] & t[23]);
  assign t[7] = t[9] | t[10];
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[23]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind216(x, y);
 input [36:0] x;
 output y;

 wire [39:0] t;
  assign t[0] = t[2] ^ t[16];
  assign t[10] = ~(t[20]);
  assign t[11] = t[13] & t[21];
  assign t[12] = ~(t[14] | t[15]);
  assign t[13] = ~(t[22] | t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = t[28] ^ x[2];
  assign t[17] = t[29] ^ x[6];
  assign t[18] = t[30] ^ x[9];
  assign t[19] = t[31] ^ x[12];
  assign t[1] = ~(t[3]);
  assign t[20] = t[32] ^ x[15];
  assign t[21] = t[33] ^ x[18];
  assign t[22] = t[34] ^ x[21];
  assign t[23] = t[35] ^ x[24];
  assign t[24] = t[36] ^ x[27];
  assign t[25] = t[37] ^ x[30];
  assign t[26] = t[38] ^ x[33];
  assign t[27] = t[39] ^ x[36];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[4] & x[5]);
  assign t[2] = t[4] | t[5];
  assign t[30] = (x[7] & x[8]);
  assign t[31] = (x[10] & x[11]);
  assign t[32] = (x[13] & x[14]);
  assign t[33] = (x[16] & x[17]);
  assign t[34] = (x[19] & x[20]);
  assign t[35] = (x[22] & x[23]);
  assign t[36] = (x[25] & x[26]);
  assign t[37] = (x[28] & x[29]);
  assign t[38] = (x[31] & x[32]);
  assign t[39] = (x[34] & x[35]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[17]);
  assign t[5] = ~(t[6] & t[18]);
  assign t[6] = t[19] & t[7];
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind217(x, y);
 input [33:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[14];
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[19] | t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = ~(t[23] & t[24]);
  assign t[14] = t[25] ^ x[2];
  assign t[15] = t[26] ^ x[5];
  assign t[16] = t[27] ^ x[9];
  assign t[17] = t[28] ^ x[12];
  assign t[18] = t[29] ^ x[15];
  assign t[19] = t[30] ^ x[18];
  assign t[1] = ~(t[3]);
  assign t[20] = t[31] ^ x[21];
  assign t[21] = t[32] ^ x[24];
  assign t[22] = t[33] ^ x[27];
  assign t[23] = t[34] ^ x[30];
  assign t[24] = t[35] ^ x[33];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[7] & x[8]);
  assign t[28] = (x[10] & x[11]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[4] & t[15]);
  assign t[30] = (x[16] & x[17]);
  assign t[31] = (x[19] & x[20]);
  assign t[32] = (x[22] & x[23]);
  assign t[33] = (x[25] & x[26]);
  assign t[34] = (x[28] & x[29]);
  assign t[35] = (x[31] & x[32]);
  assign t[3] = ~(x[6]);
  assign t[4] = t[16] & t[5];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[17]);
  assign t[9] = t[11] & t[18];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind218(x, y);
 input [30:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2] ^ t[13]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = t[23] ^ x[2];
  assign t[14] = t[24] ^ x[5];
  assign t[15] = t[25] ^ x[9];
  assign t[16] = t[26] ^ x[12];
  assign t[17] = t[27] ^ x[15];
  assign t[18] = t[28] ^ x[18];
  assign t[19] = t[29] ^ x[21];
  assign t[1] = ~(t[3]);
  assign t[20] = t[30] ^ x[24];
  assign t[21] = t[31] ^ x[27];
  assign t[22] = t[32] ^ x[30];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[7] & x[8]);
  assign t[26] = (x[10] & x[11]);
  assign t[27] = (x[13] & x[14]);
  assign t[28] = (x[16] & x[17]);
  assign t[29] = (x[19] & x[20]);
  assign t[2] = t[14] & t[4];
  assign t[30] = (x[22] & x[23]);
  assign t[31] = (x[25] & x[26]);
  assign t[32] = (x[28] & x[29]);
  assign t[3] = ~(x[6]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[15]);
  assign t[8] = t[10] & t[16];
  assign t[9] = ~(t[11] | t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind219(x, y);
 input [27:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[12] ^ t[2]);
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = t[21] ^ x[2];
  assign t[13] = t[22] ^ x[6];
  assign t[14] = t[23] ^ x[9];
  assign t[15] = t[24] ^ x[12];
  assign t[16] = t[25] ^ x[15];
  assign t[17] = t[26] ^ x[18];
  assign t[18] = t[27] ^ x[21];
  assign t[19] = t[28] ^ x[24];
  assign t[1] = ~(t[3]);
  assign t[20] = t[29] ^ x[27];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[4] & x[5]);
  assign t[23] = (x[7] & x[8]);
  assign t[24] = (x[10] & x[11]);
  assign t[25] = (x[13] & x[14]);
  assign t[26] = (x[16] & x[17]);
  assign t[27] = (x[19] & x[20]);
  assign t[28] = (x[22] & x[23]);
  assign t[29] = (x[25] & x[26]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[9] & t[14];
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind220(x, y);
 input [27:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(x[0]);
  assign t[10] = t[19] ^ x[3];
  assign t[11] = t[20] ^ x[6];
  assign t[12] = t[21] ^ x[9];
  assign t[13] = t[22] ^ x[12];
  assign t[14] = t[23] ^ x[15];
  assign t[15] = t[24] ^ x[18];
  assign t[16] = t[25] ^ x[21];
  assign t[17] = t[26] ^ x[24];
  assign t[18] = t[27] ^ x[27];
  assign t[19] = (x[1] & x[2]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[20] = (x[4] & x[5]);
  assign t[21] = (x[7] & x[8]);
  assign t[22] = (x[10] & x[11]);
  assign t[23] = (x[13] & x[14]);
  assign t[24] = (x[16] & x[17]);
  assign t[25] = (x[19] & x[20]);
  assign t[26] = (x[22] & x[23]);
  assign t[27] = (x[25] & x[26]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11] | t[12]);
  assign t[5] = ~(t[7] | t[13]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[9] = ~(t[17] & t[18]);
  assign y = t[0] & t[1];
endmodule

module R1ind221(x, y);
 input [42:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19] & t[10]);
  assign t[16] = ~(t[33] & t[20]);
  assign t[17] = ~(t[34] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[37] & t[38]);
  assign t[23] = ~(t[39] & t[40]);
  assign t[24] = ~(t[19] & t[25]);
  assign t[25] = t[26] & t[36];
  assign t[26] = ~(t[33] | t[32]);
  assign t[27] = t[41] ^ x[3];
  assign t[28] = t[42] ^ x[6];
  assign t[29] = t[43] ^ x[9];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[44] ^ x[12];
  assign t[31] = t[45] ^ x[15];
  assign t[32] = t[46] ^ x[18];
  assign t[33] = t[47] ^ x[21];
  assign t[34] = t[48] ^ x[24];
  assign t[35] = t[49] ^ x[27];
  assign t[36] = t[50] ^ x[30];
  assign t[37] = t[51] ^ x[33];
  assign t[38] = t[52] ^ x[36];
  assign t[39] = t[53] ^ x[39];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[54] ^ x[42];
  assign t[41] = (x[1] & x[2]);
  assign t[42] = (x[4] & x[5]);
  assign t[43] = (x[7] & x[8]);
  assign t[44] = (x[10] & x[11]);
  assign t[45] = (x[13] & x[14]);
  assign t[46] = (x[16] & x[17]);
  assign t[47] = (x[19] & x[20]);
  assign t[48] = (x[22] & x[23]);
  assign t[49] = (x[25] & x[26]);
  assign t[4] = ~(t[10] | t[11]);
  assign t[50] = (x[28] & x[29]);
  assign t[51] = (x[31] & x[32]);
  assign t[52] = (x[34] & x[35]);
  assign t[53] = (x[37] & x[38]);
  assign t[54] = (x[40] & x[41]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[27] & t[28]);
  assign t[7] = ~(t[29] & t[30]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[31] & t[5]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind222(x, y);
 input [42:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[30]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[31] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[32] & t[33]);
  assign t[15] = ~(t[34] & t[35]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[36] & t[7]);
  assign t[18] = ~(t[37] & t[38]);
  assign t[19] = ~(t[39] & t[40]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[41] | t[42]);
  assign t[22] = ~(t[25] | t[30]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[25] & t[28]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[25] & t[29]);
  assign t[27] = ~(t[41] & t[10]);
  assign t[28] = t[21] & t[30];
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[44] ^ x[3];
  assign t[31] = t[45] ^ x[6];
  assign t[32] = t[46] ^ x[9];
  assign t[33] = t[47] ^ x[12];
  assign t[34] = t[48] ^ x[15];
  assign t[35] = t[49] ^ x[18];
  assign t[36] = t[50] ^ x[21];
  assign t[37] = t[51] ^ x[24];
  assign t[38] = t[52] ^ x[27];
  assign t[39] = t[53] ^ x[30];
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = t[54] ^ x[33];
  assign t[41] = t[55] ^ x[36];
  assign t[42] = t[56] ^ x[39];
  assign t[43] = t[57] ^ x[42];
  assign t[44] = (x[1] & x[2]);
  assign t[45] = (x[4] & x[5]);
  assign t[46] = (x[7] & x[8]);
  assign t[47] = (x[10] & x[11]);
  assign t[48] = (x[13] & x[14]);
  assign t[49] = (x[16] & x[17]);
  assign t[4] = ~(t[10]);
  assign t[50] = (x[19] & x[20]);
  assign t[51] = (x[22] & x[23]);
  assign t[52] = (x[25] & x[26]);
  assign t[53] = (x[28] & x[29]);
  assign t[54] = (x[31] & x[32]);
  assign t[55] = (x[34] & x[35]);
  assign t[56] = (x[37] & x[38]);
  assign t[57] = (x[40] & x[41]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12] & t[13]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind223(x, y);
 input [11:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~(t[5] & t[1]);
  assign t[10] = (x[6] & x[7]);
  assign t[11] = (x[9] & x[10]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[7]);
  assign t[4] = t[8] ^ x[2];
  assign t[5] = t[9] ^ x[5];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[11];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[3] & x[4]);
  assign y = ~(t[4] | t[0]);
endmodule

module R1ind224(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind225(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind226(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind227(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind228(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[10];
  assign t[11] = t[18] ^ x[13];
  assign t[12] = t[19] ^ x[16];
  assign t[13] = t[20] ^ x[19];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[0] & x[3]);
  assign t[16] = (x[5] & x[6]);
  assign t[17] = (x[8] & x[9]);
  assign t[18] = (x[11] & x[12]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[4];
  assign t[9] = t[16] ^ x[7];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind229(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind230(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind231(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind232(x, y);
 input [12:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[14] ^ x[9];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (x[1] & x[2]);
  assign t[13] = (x[4] & x[5]);
  assign t[14] = (x[7] & x[8]);
  assign t[15] = (x[10] & x[11]);
  assign t[1] = ~(x[0]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[8] & t[7]);
  assign t[5] = ~(t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[3];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind233(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind234(x, y);
 input [17:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~(t[7] | t[2]);
  assign t[10] = t[16] ^ x[11];
  assign t[11] = t[17] ^ x[14];
  assign t[12] = t[18] ^ x[17];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[12] & x[13]);
  assign t[18] = (x[15] & x[16]);
  assign t[1] = ~(t[8]);
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = t[6] & t[10];
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = t[13] ^ x[2];
  assign t[8] = t[14] ^ x[5];
  assign t[9] = t[15] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind235(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind236(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind237(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind238(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1_ind(x, y);
 input [555:0] x;
 output [238:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[194], x[193], x[196], x[195], x[190], x[189], x[192], x[191], x[188], x[201], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[200], x[199], x[177], x[198], x[197], x[174]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[194], x[193], x[192], x[191], x[190], x[189], x[196], x[195], x[188], x[206], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[205], x[204], x[177], x[203], x[202], x[174]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[196], x[195], x[194], x[193], x[190], x[189], x[192], x[191], x[188], x[211], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[210], x[209], x[177], x[208], x[207], x[174]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[215], x[208], x[207], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[176], x[175], x[174], x[214], x[213], x[212]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[218], x[179], x[178], x[177], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[198], x[197], x[174], x[217], x[216], x[212]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[221], x[200], x[199], x[177], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[203], x[202], x[174], x[220], x[219], x[212]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[224], x[205], x[204], x[177], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[208], x[207], x[174], x[223], x[222], x[212]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[228], x[223], x[222], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[214], x[213], x[212], x[227], x[226], x[225]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[231], x[176], x[175], x[174], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[217], x[216], x[212], x[230], x[229], x[225]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[234], x[198], x[197], x[174], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[220], x[219], x[212], x[233], x[232], x[225]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[237], x[203], x[202], x[174], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[223], x[222], x[212], x[236], x[235], x[225]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[241], x[236], x[235], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[240], x[239], x[238]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[244], x[214], x[213], x[212], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[230], x[229], x[225], x[243], x[242], x[238]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[247], x[217], x[216], x[212], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[233], x[232], x[225], x[246], x[245], x[238]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[250], x[220], x[219], x[212], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[236], x[235], x[225], x[249], x[248], x[238]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[254], x[249], x[248], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[240], x[239], x[238], x[253], x[252], x[251]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[257], x[227], x[226], x[225], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[243], x[242], x[238], x[256], x[255], x[251]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[260], x[230], x[229], x[225], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[246], x[245], x[238], x[259], x[258], x[251]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[263], x[233], x[232], x[225], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[249], x[248], x[238], x[262], x[261], x[251]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[267], x[262], x[261], x[186], x[182], x[181], x[180], x[253], x[252], x[251], x[266], x[265], x[264], x[185], x[184], x[183]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[270], x[240], x[239], x[238], x[186], x[182], x[181], x[180], x[256], x[255], x[251], x[269], x[268], x[264], x[185], x[184], x[183]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[273], x[243], x[242], x[238], x[186], x[182], x[181], x[180], x[259], x[258], x[251], x[272], x[271], x[264], x[185], x[184], x[183]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[276], x[246], x[245], x[238], x[186], x[182], x[181], x[180], x[262], x[261], x[251], x[275], x[274], x[264], x[185], x[184], x[183]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[280], x[275], x[274], x[186], x[182], x[181], x[180], x[266], x[265], x[264], x[279], x[278], x[277], x[185], x[184], x[183]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[283], x[253], x[252], x[251], x[186], x[182], x[181], x[180], x[269], x[268], x[264], x[282], x[281], x[277], x[185], x[184], x[183]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[286], x[256], x[255], x[251], x[186], x[182], x[181], x[180], x[272], x[271], x[264], x[285], x[284], x[277], x[185], x[184], x[183]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[289], x[259], x[258], x[251], x[186], x[182], x[181], x[180], x[275], x[274], x[264], x[288], x[287], x[277], x[185], x[184], x[183]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[296], x[288], x[287], x[186], x[295], x[294], x[293], x[279], x[278], x[277], x[292], x[291], x[290], x[185], x[184], x[183]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[299], x[266], x[265], x[264], x[186], x[295], x[294], x[293], x[282], x[281], x[277], x[298], x[297], x[290], x[185], x[184], x[183]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[302], x[269], x[268], x[264], x[186], x[295], x[294], x[293], x[285], x[284], x[277], x[301], x[300], x[290], x[185], x[184], x[183]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[305], x[272], x[271], x[264], x[186], x[295], x[294], x[293], x[288], x[287], x[277], x[304], x[303], x[290], x[185], x[184], x[183]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[312], x[304], x[303], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[292], x[291], x[290], x[308], x[307], x[306]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[315], x[279], x[278], x[277], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[298], x[297], x[290], x[314], x[313], x[306]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[318], x[282], x[281], x[277], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[301], x[300], x[290], x[317], x[316], x[306]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[321], x[285], x[284], x[277], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[304], x[303], x[290], x[320], x[319], x[306]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[325], x[320], x[319], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[308], x[307], x[306], x[324], x[323], x[322]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[328], x[292], x[291], x[290], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[314], x[313], x[306], x[327], x[326], x[322]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[331], x[298], x[297], x[290], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[317], x[316], x[306], x[330], x[329], x[322]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[334], x[301], x[300], x[290], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[320], x[319], x[306], x[333], x[332], x[322]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[338], x[333], x[332], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[324], x[323], x[322], x[337], x[336], x[335]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[341], x[308], x[307], x[306], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[327], x[326], x[322], x[340], x[339], x[335]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[344], x[314], x[313], x[306], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[330], x[329], x[322], x[343], x[342], x[335]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[347], x[317], x[316], x[306], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[333], x[332], x[322], x[346], x[345], x[335]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[351], x[346], x[345], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[337], x[336], x[335], x[350], x[349], x[348]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[354], x[324], x[323], x[322], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[340], x[339], x[335], x[353], x[352], x[348]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[357], x[327], x[326], x[322], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[343], x[342], x[335], x[356], x[355], x[348]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[360], x[330], x[329], x[322], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[346], x[345], x[335], x[359], x[358], x[348]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[364], x[359], x[358], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[350], x[349], x[348], x[363], x[362], x[361]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[367], x[337], x[336], x[335], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[353], x[352], x[348], x[366], x[365], x[361]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[370], x[340], x[339], x[335], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[356], x[355], x[348], x[369], x[368], x[361]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[373], x[343], x[342], x[335], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[359], x[358], x[348], x[372], x[371], x[361]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[377], x[372], x[371], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[363], x[362], x[361], x[376], x[375], x[374]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[380], x[350], x[349], x[348], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[366], x[365], x[361], x[379], x[378], x[374]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[383], x[353], x[352], x[348], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[369], x[368], x[361], x[382], x[381], x[374]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[386], x[356], x[355], x[348], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[372], x[371], x[361], x[385], x[384], x[374]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[393], x[385], x[384], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[376], x[375], x[374], x[389], x[388], x[387]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[396], x[363], x[362], x[361], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[379], x[378], x[374], x[395], x[394], x[387]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[399], x[366], x[365], x[361], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[382], x[381], x[374], x[398], x[397], x[387]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[402], x[369], x[368], x[361], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[385], x[384], x[374], x[401], x[400], x[387]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[401], x[400], x[409], x[408], x[407], x[406], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[389], x[388], x[387], x[405], x[404], x[403]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[376], x[375], x[374], x[415], x[414], x[413], x[412], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[395], x[394], x[387], x[411], x[410], x[403]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[379], x[378], x[374], x[421], x[420], x[419], x[418], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[398], x[397], x[387], x[417], x[416], x[403]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[382], x[381], x[374], x[427], x[426], x[425], x[424], x[186], x[311], x[310], x[309], x[392], x[391], x[390], x[401], x[400], x[387], x[423], x[422], x[403]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[431], x[423], x[422], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[405], x[404], x[403], x[430], x[429], x[428]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[434], x[389], x[388], x[387], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[411], x[410], x[403], x[433], x[432], x[428]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[437], x[395], x[394], x[387], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[417], x[416], x[403], x[436], x[435], x[428]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[398], x[397], x[387], x[443], x[442], x[441], x[440], x[186], x[311], x[310], x[309], x[295], x[294], x[293], x[423], x[422], x[403], x[439], x[438], x[428]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[447], x[439], x[438], x[186], x[311], x[310], x[309], x[182], x[181], x[180], x[430], x[429], x[428], x[446], x[445], x[444]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[450], x[405], x[404], x[403], x[186], x[311], x[310], x[309], x[182], x[181], x[180], x[433], x[432], x[428], x[449], x[448], x[444]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[453], x[411], x[410], x[403], x[186], x[311], x[310], x[309], x[182], x[181], x[180], x[436], x[435], x[428], x[452], x[451], x[444]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[456], x[417], x[416], x[403], x[186], x[311], x[310], x[309], x[182], x[181], x[180], x[439], x[438], x[428], x[455], x[454], x[444]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[460], x[455], x[454], x[186], x[295], x[294], x[293], x[446], x[445], x[444], x[459], x[458], x[457], x[311], x[310], x[309]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[463], x[430], x[429], x[428], x[186], x[295], x[294], x[293], x[449], x[448], x[444], x[462], x[461], x[457], x[311], x[310], x[309]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[466], x[433], x[432], x[428], x[186], x[295], x[294], x[293], x[452], x[451], x[444], x[465], x[464], x[457], x[311], x[310], x[309]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[469], x[436], x[435], x[428], x[186], x[295], x[294], x[293], x[455], x[454], x[444], x[468], x[467], x[457], x[311], x[310], x[309]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[470], x[468], x[467], x[186], x[182], x[181], x[180], x[459], x[458], x[457], x[179], x[178], x[177], x[311], x[310], x[309]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[471], x[446], x[445], x[444], x[186], x[182], x[181], x[180], x[462], x[461], x[457], x[200], x[199], x[177], x[311], x[310], x[309]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[472], x[449], x[448], x[444], x[186], x[182], x[181], x[180], x[465], x[464], x[457], x[205], x[204], x[177], x[311], x[310], x[309]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[473], x[452], x[451], x[444], x[186], x[182], x[181], x[180], x[468], x[467], x[457], x[210], x[209], x[177], x[311], x[310], x[309]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[186], x[480], x[113], x[112], x[111], x[479], x[478], x[477], x[476], x[475], x[474], x[146], x[145], x[138], x[137], x[136], x[129]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[186], x[481], x[122], x[121], x[120], x[479], x[478], x[477], x[476], x[475], x[474], x[144], x[143], x[138], x[135], x[134], x[129]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[482], x[131], x[130], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[142], x[141], x[138], x[133], x[132], x[129]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[186], x[483], x[479], x[478], x[477], x[476], x[475], x[474], x[140], x[139], x[138], x[131], x[130], x[129]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[484], x[77], x[76], x[75], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[137], x[136], x[129], x[128], x[127], x[120]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[485], x[86], x[85], x[84], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[135], x[134], x[129], x[126], x[125], x[120]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[486], x[95], x[94], x[93], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[133], x[132], x[129], x[124], x[123], x[120]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[487], x[104], x[103], x[102], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[131], x[130], x[129], x[122], x[121], x[120]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[488], x[41], x[40], x[39], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[128], x[127], x[120], x[119], x[118], x[111]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[489], x[50], x[49], x[48], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[126], x[125], x[120], x[117], x[116], x[111]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[490], x[59], x[58], x[57], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[124], x[123], x[120], x[115], x[114], x[111]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[491], x[68], x[67], x[66], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[122], x[121], x[120], x[113], x[112], x[111]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[186], x[492], x[11], x[10], x[3], x[479], x[478], x[477], x[476], x[475], x[474], x[119], x[118], x[111], x[110], x[109], x[102]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[186], x[493], x[14], x[13], x[12], x[479], x[478], x[477], x[476], x[475], x[474], x[117], x[116], x[111], x[108], x[107], x[102]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[186], x[494], x[23], x[22], x[21], x[479], x[478], x[477], x[476], x[475], x[474], x[115], x[114], x[111], x[106], x[105], x[102]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[495], x[32], x[31], x[30], x[186], x[479], x[478], x[477], x[476], x[475], x[474], x[113], x[112], x[111], x[104], x[103], x[102]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[496], x[115], x[114], x[111], x[186], x[476], x[475], x[474], x[110], x[109], x[102], x[101], x[100], x[93], x[479], x[478], x[477]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[497], x[124], x[123], x[120], x[186], x[476], x[475], x[474], x[108], x[107], x[102], x[99], x[98], x[93], x[479], x[478], x[477]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[186], x[498], x[133], x[132], x[129], x[476], x[475], x[474], x[106], x[105], x[102], x[97], x[96], x[93], x[479], x[478], x[477]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[186], x[499], x[142], x[141], x[138], x[476], x[475], x[474], x[104], x[103], x[102], x[95], x[94], x[93], x[479], x[478], x[477]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[500], x[79], x[78], x[75], x[186], x[476], x[475], x[474], x[101], x[100], x[93], x[92], x[91], x[84], x[479], x[478], x[477]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[186], x[501], x[88], x[87], x[476], x[475], x[474], x[99], x[98], x[93], x[90], x[89], x[84], x[479], x[478], x[477]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[186], x[502], x[476], x[475], x[474], x[97], x[96], x[93], x[88], x[87], x[84], x[479], x[478], x[477]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[503], x[106], x[105], x[102], x[186], x[476], x[475], x[474], x[95], x[94], x[93], x[86], x[85], x[84], x[479], x[478], x[477]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[186], x[504], x[43], x[42], x[39], x[476], x[475], x[474], x[92], x[91], x[84], x[83], x[82], x[75], x[479], x[478], x[477]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[186], x[505], x[52], x[51], x[48], x[476], x[475], x[474], x[90], x[89], x[84], x[81], x[80], x[75], x[479], x[478], x[477]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[186], x[506], x[61], x[60], x[57], x[476], x[475], x[474], x[88], x[87], x[84], x[79], x[78], x[75], x[479], x[478], x[477]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[507], x[70], x[69], x[66], x[186], x[476], x[475], x[474], x[86], x[85], x[84], x[77], x[76], x[75], x[479], x[478], x[477]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[186], x[511], x[9], x[8], x[3], x[479], x[478], x[477], x[510], x[509], x[508], x[83], x[82], x[75], x[74], x[73], x[66]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[186], x[512], x[16], x[15], x[12], x[479], x[478], x[477], x[510], x[509], x[508], x[81], x[80], x[75], x[72], x[71], x[66]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[186], x[513], x[25], x[24], x[21], x[479], x[478], x[477], x[510], x[509], x[508], x[79], x[78], x[75], x[70], x[69], x[66]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[186], x[514], x[34], x[33], x[30], x[479], x[478], x[477], x[510], x[509], x[508], x[77], x[76], x[75], x[68], x[67], x[66]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[186], x[515], x[117], x[116], x[111], x[479], x[478], x[477], x[510], x[509], x[508], x[74], x[73], x[66], x[65], x[64], x[57]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[186], x[516], x[126], x[125], x[120], x[479], x[478], x[477], x[510], x[509], x[508], x[72], x[71], x[66], x[63], x[62], x[57]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[186], x[517], x[135], x[134], x[129], x[479], x[478], x[477], x[510], x[509], x[508], x[70], x[69], x[66], x[61], x[60], x[57]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[186], x[518], x[144], x[143], x[138], x[479], x[478], x[477], x[510], x[509], x[508], x[68], x[67], x[66], x[59], x[58], x[57]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[186], x[519], x[81], x[80], x[75], x[479], x[478], x[477], x[510], x[509], x[508], x[65], x[64], x[57], x[56], x[55], x[48]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[186], x[520], x[90], x[89], x[84], x[479], x[478], x[477], x[510], x[509], x[508], x[63], x[62], x[57], x[54], x[53], x[48]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[186], x[521], x[99], x[98], x[93], x[479], x[478], x[477], x[510], x[509], x[508], x[61], x[60], x[57], x[52], x[51], x[48]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[186], x[522], x[108], x[107], x[102], x[479], x[478], x[477], x[510], x[509], x[508], x[59], x[58], x[57], x[50], x[49], x[48]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[186], x[523], x[45], x[44], x[479], x[478], x[477], x[510], x[509], x[508], x[56], x[55], x[48], x[47], x[46], x[39]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[186], x[524], x[479], x[478], x[477], x[510], x[509], x[508], x[54], x[53], x[48], x[45], x[44], x[39]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[186], x[525], x[63], x[62], x[57], x[479], x[478], x[477], x[510], x[509], x[508], x[52], x[51], x[48], x[43], x[42], x[39]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[186], x[526], x[72], x[71], x[66], x[479], x[478], x[477], x[510], x[509], x[508], x[50], x[49], x[48], x[41], x[40], x[39]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[186], x[527], x[7], x[6], x[3], x[510], x[509], x[508], x[47], x[46], x[39], x[38], x[37], x[30], x[479], x[478], x[477]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[186], x[528], x[18], x[17], x[12], x[510], x[509], x[508], x[45], x[44], x[39], x[36], x[35], x[30], x[479], x[478], x[477]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[186], x[529], x[27], x[26], x[21], x[510], x[509], x[508], x[43], x[42], x[39], x[34], x[33], x[30], x[479], x[478], x[477]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[186], x[530], x[36], x[35], x[510], x[509], x[508], x[41], x[40], x[39], x[32], x[31], x[30], x[479], x[478], x[477]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[186], x[531], x[119], x[118], x[111], x[479], x[478], x[477], x[510], x[509], x[508], x[38], x[37], x[30], x[29], x[28], x[21]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[186], x[532], x[128], x[127], x[120], x[479], x[478], x[477], x[510], x[509], x[508], x[36], x[35], x[30], x[27], x[26], x[21]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[186], x[533], x[137], x[136], x[129], x[479], x[478], x[477], x[510], x[509], x[508], x[34], x[33], x[30], x[25], x[24], x[21]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[186], x[534], x[146], x[145], x[138], x[479], x[478], x[477], x[510], x[509], x[508], x[32], x[31], x[30], x[23], x[22], x[21]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[186], x[535], x[83], x[82], x[75], x[479], x[478], x[477], x[510], x[509], x[508], x[29], x[28], x[21], x[20], x[19], x[12]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[186], x[536], x[92], x[91], x[84], x[479], x[478], x[477], x[510], x[509], x[508], x[27], x[26], x[21], x[18], x[17], x[12]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[186], x[537], x[101], x[100], x[93], x[479], x[478], x[477], x[510], x[509], x[508], x[25], x[24], x[21], x[16], x[15], x[12]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[186], x[538], x[110], x[109], x[102], x[479], x[478], x[477], x[510], x[509], x[508], x[23], x[22], x[21], x[14], x[13], x[12]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[186], x[539], x[47], x[46], x[39], x[479], x[478], x[477], x[392], x[391], x[390], x[20], x[19], x[12], x[5], x[4], x[3]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[186], x[540], x[56], x[55], x[48], x[479], x[478], x[477], x[392], x[391], x[390], x[18], x[17], x[12], x[7], x[6], x[3]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[186], x[541], x[65], x[64], x[57], x[479], x[478], x[477], x[392], x[391], x[390], x[16], x[15], x[12], x[9], x[8], x[3]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[186], x[542], x[74], x[73], x[66], x[479], x[478], x[477], x[392], x[391], x[390], x[14], x[13], x[12], x[11], x[10], x[3]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[196], x[195], x[186], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[146], x[145], x[138], x[179], x[178], x[177], x[543], x[149], x[148], x[147], x[392], x[391], x[390], x[5], x[4], x[3], x[479], x[478], x[477]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[194], x[193], x[196], x[195], x[190], x[189], x[192], x[191], x[188], x[186], x[144], x[143], x[138], x[200], x[199], x[177], x[544], x[20], x[19], x[12], x[149], x[148], x[147], x[392], x[391], x[390], x[7], x[6], x[3], x[479], x[478], x[477]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[194], x[193], x[192], x[191], x[190], x[189], x[196], x[195], x[188], x[186], x[142], x[141], x[138], x[205], x[204], x[177], x[545], x[29], x[28], x[21], x[149], x[148], x[147], x[392], x[391], x[390], x[9], x[8], x[3], x[479], x[478], x[477]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[196], x[195], x[194], x[193], x[190], x[189], x[186], x[192], x[191], x[188], x[140], x[139], x[138], x[210], x[209], x[177], x[546], x[38], x[37], x[30], x[149], x[148], x[147], x[392], x[391], x[390], x[11], x[10], x[3], x[479], x[478], x[477]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[186]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[149], x[148], x[147], x[170], x[169], x[168], x[173], x[172], x[171], x[164], x[163], x[162], x[392], x[391], x[390], x[167], x[166], x[165]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[149], x[148], x[147], x[170], x[169], x[168], x[173], x[172], x[171], x[392], x[391], x[390], x[164], x[163], x[162]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[149], x[148], x[147], x[170], x[169], x[168], x[392], x[391], x[390], x[173], x[172], x[171]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[149], x[148], x[147], x[170], x[169], x[168], x[392], x[391], x[390]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[443], x[442], x[441], x[409], x[408], x[407], x[415], x[414], x[413], x[421], x[420], x[419], x[186], x[427], x[426], x[425]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[443], x[442], x[441], x[409], x[408], x[407], x[415], x[414], x[413], x[186], x[421], x[420], x[419]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[443], x[442], x[441], x[186], x[409], x[408], x[407], x[415], x[414], x[413]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[186], x[443], x[442], x[441], x[409], x[408], x[407]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[186], x[443], x[442], x[441]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[186]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[158], x[157], x[156], x[161], x[160], x[159], x[149], x[148], x[147], x[152], x[151], x[150], x[155], x[154], x[153], x[443], x[442], x[441], x[427], x[426], x[425], x[415], x[414], x[413], x[421], x[420], x[419], x[409], x[408], x[407], x[186]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[161], x[160], x[159], x[155], x[154], x[153], x[152], x[151], x[150], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[443], x[442], x[441], x[427], x[426], x[425], x[415], x[414], x[413], x[421], x[420], x[419], x[409], x[408], x[407], x[149], x[148], x[147], x[158], x[157], x[156], x[186]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[158], x[157], x[156], x[161], x[160], x[159], x[155], x[154], x[153], x[152], x[151], x[150]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[549], x[548], x[547]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[552], x[551], x[550]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[161], x[160], x[159], x[152], x[151], x[150], x[144], x[143], x[138], x[200], x[199], x[177], x[459], x[458], x[457]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[161], x[160], x[159], x[152], x[151], x[150], x[140], x[139], x[138], x[210], x[209], x[177], x[465], x[464], x[457]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[161], x[160], x[159], x[152], x[151], x[150], x[146], x[145], x[138], x[179], x[178], x[210], x[209], x[177]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[161], x[160], x[159], x[152], x[151], x[150], x[142], x[141], x[138], x[205], x[204], x[177], x[462], x[461], x[457]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[549], x[548], x[547]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[552], x[551], x[550]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[161], x[160], x[159], x[152], x[151], x[150], x[186]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[555], x[554], x[553]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[161], x[160], x[159], x[392], x[391], x[390], x[149], x[148], x[147]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[555], x[554], x[553]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[392], x[391], x[390]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[479], x[478], x[477]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[392], x[391], x[390]}), .y(y[238]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[5];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[29] ^ x[8];
  assign t[21] = t[30] ^ x[11];
  assign t[22] = t[31] ^ x[14];
  assign t[23] = t[32] ^ x[17];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[23];
  assign t[26] = t[35] ^ x[26];
  assign t[27] = (~t[36] & t[37]);
  assign t[28] = (~t[38] & t[39]);
  assign t[29] = (~t[40] & t[41]);
  assign t[2] = ~(t[9] & t[5]);
  assign t[30] = (~t[42] & t[43]);
  assign t[31] = (~t[44] & t[45]);
  assign t[32] = (~t[46] & t[47]);
  assign t[33] = (~t[48] & t[49]);
  assign t[34] = (~t[50] & t[51]);
  assign t[35] = (~t[52] & t[53]);
  assign t[36] = t[54] ^ x[1];
  assign t[37] = t[55] ^ x[2];
  assign t[38] = t[56] ^ x[4];
  assign t[39] = t[57] ^ x[5];
  assign t[3] = ~(t[10] | t[11]);
  assign t[40] = t[58] ^ x[7];
  assign t[41] = t[59] ^ x[8];
  assign t[42] = t[60] ^ x[10];
  assign t[43] = t[61] ^ x[11];
  assign t[44] = t[62] ^ x[13];
  assign t[45] = t[63] ^ x[14];
  assign t[46] = t[64] ^ x[16];
  assign t[47] = t[65] ^ x[17];
  assign t[48] = t[66] ^ x[19];
  assign t[49] = t[67] ^ x[20];
  assign t[4] = ~(t[6] | t[12]);
  assign t[50] = t[68] ^ x[22];
  assign t[51] = t[69] ^ x[23];
  assign t[52] = t[70] ^ x[25];
  assign t[53] = t[71] ^ x[26];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13]);
  assign t[70] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[24]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[8] = ~(t[16] & t[17]);
  assign t[9] = (t[18]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[5];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[29] ^ x[8];
  assign t[21] = t[30] ^ x[11];
  assign t[22] = t[31] ^ x[14];
  assign t[23] = t[32] ^ x[17];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[23];
  assign t[26] = t[35] ^ x[26];
  assign t[27] = (~t[36] & t[37]);
  assign t[28] = (~t[38] & t[39]);
  assign t[29] = (~t[40] & t[41]);
  assign t[2] = ~(t[9] & t[5]);
  assign t[30] = (~t[42] & t[43]);
  assign t[31] = (~t[44] & t[45]);
  assign t[32] = (~t[46] & t[47]);
  assign t[33] = (~t[48] & t[49]);
  assign t[34] = (~t[50] & t[51]);
  assign t[35] = (~t[52] & t[53]);
  assign t[36] = t[54] ^ x[1];
  assign t[37] = t[55] ^ x[2];
  assign t[38] = t[56] ^ x[4];
  assign t[39] = t[57] ^ x[5];
  assign t[3] = ~(t[10] | t[11]);
  assign t[40] = t[58] ^ x[7];
  assign t[41] = t[59] ^ x[8];
  assign t[42] = t[60] ^ x[10];
  assign t[43] = t[61] ^ x[11];
  assign t[44] = t[62] ^ x[13];
  assign t[45] = t[63] ^ x[14];
  assign t[46] = t[64] ^ x[16];
  assign t[47] = t[65] ^ x[17];
  assign t[48] = t[66] ^ x[19];
  assign t[49] = t[67] ^ x[20];
  assign t[4] = ~(t[6] | t[12]);
  assign t[50] = t[68] ^ x[22];
  assign t[51] = t[69] ^ x[23];
  assign t[52] = t[70] ^ x[25];
  assign t[53] = t[71] ^ x[26];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13]);
  assign t[70] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[24]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[8] = ~(t[16] & t[17]);
  assign t[9] = (t[18]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = (~t[47] & t[48]);
  assign t[34] = (~t[49] & t[50]);
  assign t[35] = t[51] ^ x[2];
  assign t[36] = t[52] ^ x[3];
  assign t[37] = t[53] ^ x[5];
  assign t[38] = t[54] ^ x[6];
  assign t[39] = t[55] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[9];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[12];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[15];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[18];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[21];
  assign t[49] = t[65] ^ x[23];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[24];
  assign t[51] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[1]);
  assign t[53] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[4]);
  assign t[55] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[7]);
  assign t[57] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[10]);
  assign t[59] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[16]);
  assign t[63] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[19]);
  assign t[65] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = (~t[47] & t[48]);
  assign t[34] = (~t[49] & t[50]);
  assign t[35] = t[51] ^ x[2];
  assign t[36] = t[52] ^ x[3];
  assign t[37] = t[53] ^ x[5];
  assign t[38] = t[54] ^ x[6];
  assign t[39] = t[55] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[9];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[12];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[15];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[18];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[21];
  assign t[49] = t[65] ^ x[23];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[24];
  assign t[51] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[1]);
  assign t[53] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[4]);
  assign t[55] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[7]);
  assign t[57] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[10]);
  assign t[59] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[16]);
  assign t[63] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[19]);
  assign t[65] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [42:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[4]);
  assign t[102] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[103] = (x[7]);
  assign t[104] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[10]);
  assign t[106] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[107] = (x[13]);
  assign t[108] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[16]);
  assign t[10] = ~(t[32] & t[6]);
  assign t[110] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[111] = (x[19]);
  assign t[112] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[113] = (x[22]);
  assign t[114] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[115] = (x[25]);
  assign t[116] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[28]);
  assign t[118] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[31]);
  assign t[11] = ~(t[33]);
  assign t[120] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[34]);
  assign t[122] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[37]);
  assign t[124] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[40]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[34] & t[21]);
  assign t[18] = ~(t[35] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[38] & t[39]);
  assign t[24] = ~(t[40] & t[41]);
  assign t[25] = ~(t[20] & t[26]);
  assign t[26] = t[27] & t[37];
  assign t[27] = ~(t[34] | t[33]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = t[56] ^ x[3];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[12];
  assign t[46] = t[60] ^ x[15];
  assign t[47] = t[61] ^ x[18];
  assign t[48] = t[62] ^ x[21];
  assign t[49] = t[63] ^ x[24];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[64] ^ x[27];
  assign t[51] = t[65] ^ x[30];
  assign t[52] = t[66] ^ x[33];
  assign t[53] = t[67] ^ x[36];
  assign t[54] = t[68] ^ x[39];
  assign t[55] = t[69] ^ x[42];
  assign t[56] = (~t[70] & t[71]);
  assign t[57] = (~t[72] & t[73]);
  assign t[58] = (~t[74] & t[75]);
  assign t[59] = (~t[76] & t[77]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (~t[78] & t[79]);
  assign t[61] = (~t[80] & t[81]);
  assign t[62] = (~t[82] & t[83]);
  assign t[63] = (~t[84] & t[85]);
  assign t[64] = (~t[86] & t[87]);
  assign t[65] = (~t[88] & t[89]);
  assign t[66] = (~t[90] & t[91]);
  assign t[67] = (~t[92] & t[93]);
  assign t[68] = (~t[94] & t[95]);
  assign t[69] = (~t[96] & t[97]);
  assign t[6] = ~(x[0]);
  assign t[70] = t[98] ^ x[2];
  assign t[71] = t[99] ^ x[3];
  assign t[72] = t[100] ^ x[5];
  assign t[73] = t[101] ^ x[6];
  assign t[74] = t[102] ^ x[8];
  assign t[75] = t[103] ^ x[9];
  assign t[76] = t[104] ^ x[11];
  assign t[77] = t[105] ^ x[12];
  assign t[78] = t[106] ^ x[14];
  assign t[79] = t[107] ^ x[15];
  assign t[7] = ~(t[28] & t[29]);
  assign t[80] = t[108] ^ x[17];
  assign t[81] = t[109] ^ x[18];
  assign t[82] = t[110] ^ x[20];
  assign t[83] = t[111] ^ x[21];
  assign t[84] = t[112] ^ x[23];
  assign t[85] = t[113] ^ x[24];
  assign t[86] = t[114] ^ x[26];
  assign t[87] = t[115] ^ x[27];
  assign t[88] = t[116] ^ x[29];
  assign t[89] = t[117] ^ x[30];
  assign t[8] = ~(t[30] & t[31]);
  assign t[90] = t[118] ^ x[32];
  assign t[91] = t[119] ^ x[33];
  assign t[92] = t[120] ^ x[35];
  assign t[93] = t[121] ^ x[36];
  assign t[94] = t[122] ^ x[38];
  assign t[95] = t[123] ^ x[39];
  assign t[96] = t[124] ^ x[41];
  assign t[97] = t[125] ^ x[42];
  assign t[98] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[1]);
  assign t[9] = ~(t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [42:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[4]);
  assign t[102] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[103] = (x[7]);
  assign t[104] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[10]);
  assign t[106] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[107] = (x[13]);
  assign t[108] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[16]);
  assign t[10] = ~(t[32] & t[6]);
  assign t[110] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[111] = (x[19]);
  assign t[112] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[113] = (x[22]);
  assign t[114] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[115] = (x[25]);
  assign t[116] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[28]);
  assign t[118] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[31]);
  assign t[11] = ~(t[33]);
  assign t[120] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[34]);
  assign t[122] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[37]);
  assign t[124] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[40]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[34] & t[21]);
  assign t[18] = ~(t[35] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[38] & t[39]);
  assign t[24] = ~(t[40] & t[41]);
  assign t[25] = ~(t[20] & t[26]);
  assign t[26] = t[27] & t[37];
  assign t[27] = ~(t[34] | t[33]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = t[56] ^ x[3];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[12];
  assign t[46] = t[60] ^ x[15];
  assign t[47] = t[61] ^ x[18];
  assign t[48] = t[62] ^ x[21];
  assign t[49] = t[63] ^ x[24];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[64] ^ x[27];
  assign t[51] = t[65] ^ x[30];
  assign t[52] = t[66] ^ x[33];
  assign t[53] = t[67] ^ x[36];
  assign t[54] = t[68] ^ x[39];
  assign t[55] = t[69] ^ x[42];
  assign t[56] = (~t[70] & t[71]);
  assign t[57] = (~t[72] & t[73]);
  assign t[58] = (~t[74] & t[75]);
  assign t[59] = (~t[76] & t[77]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (~t[78] & t[79]);
  assign t[61] = (~t[80] & t[81]);
  assign t[62] = (~t[82] & t[83]);
  assign t[63] = (~t[84] & t[85]);
  assign t[64] = (~t[86] & t[87]);
  assign t[65] = (~t[88] & t[89]);
  assign t[66] = (~t[90] & t[91]);
  assign t[67] = (~t[92] & t[93]);
  assign t[68] = (~t[94] & t[95]);
  assign t[69] = (~t[96] & t[97]);
  assign t[6] = ~(x[0]);
  assign t[70] = t[98] ^ x[2];
  assign t[71] = t[99] ^ x[3];
  assign t[72] = t[100] ^ x[5];
  assign t[73] = t[101] ^ x[6];
  assign t[74] = t[102] ^ x[8];
  assign t[75] = t[103] ^ x[9];
  assign t[76] = t[104] ^ x[11];
  assign t[77] = t[105] ^ x[12];
  assign t[78] = t[106] ^ x[14];
  assign t[79] = t[107] ^ x[15];
  assign t[7] = ~(t[28] & t[29]);
  assign t[80] = t[108] ^ x[17];
  assign t[81] = t[109] ^ x[18];
  assign t[82] = t[110] ^ x[20];
  assign t[83] = t[111] ^ x[21];
  assign t[84] = t[112] ^ x[23];
  assign t[85] = t[113] ^ x[24];
  assign t[86] = t[114] ^ x[26];
  assign t[87] = t[115] ^ x[27];
  assign t[88] = t[116] ^ x[29];
  assign t[89] = t[117] ^ x[30];
  assign t[8] = ~(t[30] & t[31]);
  assign t[90] = t[118] ^ x[32];
  assign t[91] = t[119] ^ x[33];
  assign t[92] = t[120] ^ x[35];
  assign t[93] = t[121] ^ x[36];
  assign t[94] = t[122] ^ x[38];
  assign t[95] = t[123] ^ x[39];
  assign t[96] = t[124] ^ x[41];
  assign t[97] = t[125] ^ x[42];
  assign t[98] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[1]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [27:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[18] & t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(x[0]);
  assign t[20] = t[29] ^ x[3];
  assign t[21] = t[30] ^ x[6];
  assign t[22] = t[31] ^ x[9];
  assign t[23] = t[32] ^ x[12];
  assign t[24] = t[33] ^ x[15];
  assign t[25] = t[34] ^ x[18];
  assign t[26] = t[35] ^ x[21];
  assign t[27] = t[36] ^ x[24];
  assign t[28] = t[37] ^ x[27];
  assign t[29] = (~t[38] & t[39]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (~t[40] & t[41]);
  assign t[31] = (~t[42] & t[43]);
  assign t[32] = (~t[44] & t[45]);
  assign t[33] = (~t[46] & t[47]);
  assign t[34] = (~t[48] & t[49]);
  assign t[35] = (~t[50] & t[51]);
  assign t[36] = (~t[52] & t[53]);
  assign t[37] = (~t[54] & t[55]);
  assign t[38] = t[56] ^ x[2];
  assign t[39] = t[57] ^ x[3];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[58] ^ x[5];
  assign t[41] = t[59] ^ x[6];
  assign t[42] = t[60] ^ x[8];
  assign t[43] = t[61] ^ x[9];
  assign t[44] = t[62] ^ x[11];
  assign t[45] = t[63] ^ x[12];
  assign t[46] = t[64] ^ x[14];
  assign t[47] = t[65] ^ x[15];
  assign t[48] = t[66] ^ x[17];
  assign t[49] = t[67] ^ x[18];
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = t[68] ^ x[20];
  assign t[51] = t[69] ^ x[21];
  assign t[52] = t[70] ^ x[23];
  assign t[53] = t[71] ^ x[24];
  assign t[54] = t[72] ^ x[26];
  assign t[55] = t[73] ^ x[27];
  assign t[56] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[1]);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[12] | t[13]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[68] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[8] | t[14]);
  assign t[70] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[22]);
  assign t[72] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[25]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [27:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[18] & t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(x[0]);
  assign t[20] = t[29] ^ x[3];
  assign t[21] = t[30] ^ x[6];
  assign t[22] = t[31] ^ x[9];
  assign t[23] = t[32] ^ x[12];
  assign t[24] = t[33] ^ x[15];
  assign t[25] = t[34] ^ x[18];
  assign t[26] = t[35] ^ x[21];
  assign t[27] = t[36] ^ x[24];
  assign t[28] = t[37] ^ x[27];
  assign t[29] = (~t[38] & t[39]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (~t[40] & t[41]);
  assign t[31] = (~t[42] & t[43]);
  assign t[32] = (~t[44] & t[45]);
  assign t[33] = (~t[46] & t[47]);
  assign t[34] = (~t[48] & t[49]);
  assign t[35] = (~t[50] & t[51]);
  assign t[36] = (~t[52] & t[53]);
  assign t[37] = (~t[54] & t[55]);
  assign t[38] = t[56] ^ x[2];
  assign t[39] = t[57] ^ x[3];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[58] ^ x[5];
  assign t[41] = t[59] ^ x[6];
  assign t[42] = t[60] ^ x[8];
  assign t[43] = t[61] ^ x[9];
  assign t[44] = t[62] ^ x[11];
  assign t[45] = t[63] ^ x[12];
  assign t[46] = t[64] ^ x[14];
  assign t[47] = t[65] ^ x[15];
  assign t[48] = t[66] ^ x[17];
  assign t[49] = t[67] ^ x[18];
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = t[68] ^ x[20];
  assign t[51] = t[69] ^ x[21];
  assign t[52] = t[70] ^ x[23];
  assign t[53] = t[71] ^ x[24];
  assign t[54] = t[72] ^ x[26];
  assign t[55] = t[73] ^ x[27];
  assign t[56] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[1]);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[12] | t[13]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[68] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[8] | t[14]);
  assign t[70] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[22]);
  assign t[72] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[25]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [42:0] x;
 output y;

 wire [128:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[128] ^ x[42];
  assign t[101] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[1]);
  assign t[103] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[4]);
  assign t[105] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[7]);
  assign t[107] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[10]);
  assign t[109] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[13]);
  assign t[111] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[16]);
  assign t[113] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[19]);
  assign t[115] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[22]);
  assign t[117] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[25]);
  assign t[119] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[31]);
  assign t[120] = (x[28]);
  assign t[121] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[31]);
  assign t[123] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[34]);
  assign t[125] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[37]);
  assign t[127] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[40]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[32] | t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[33] & t[34]);
  assign t[16] = ~(t[35] & t[36]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[37] & t[8]);
  assign t[19] = ~(t[38] & t[39]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[40] & t[41]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[26] | t[31]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[26] & t[29]);
  assign t[26] = ~(t[44]);
  assign t[27] = ~(t[26] & t[30]);
  assign t[28] = ~(t[42] & t[11]);
  assign t[29] = t[22] & t[31];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[43]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = t[59] ^ x[3];
  assign t[46] = t[60] ^ x[6];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[15];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[21];
  assign t[52] = t[66] ^ x[24];
  assign t[53] = t[67] ^ x[27];
  assign t[54] = t[68] ^ x[30];
  assign t[55] = t[69] ^ x[33];
  assign t[56] = t[70] ^ x[36];
  assign t[57] = t[71] ^ x[39];
  assign t[58] = t[72] ^ x[42];
  assign t[59] = (~t[73] & t[74]);
  assign t[5] = ~(t[11]);
  assign t[60] = (~t[75] & t[76]);
  assign t[61] = (~t[77] & t[78]);
  assign t[62] = (~t[79] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[87] & t[88]);
  assign t[67] = (~t[89] & t[90]);
  assign t[68] = (~t[91] & t[92]);
  assign t[69] = (~t[93] & t[94]);
  assign t[6] = ~(t[12]);
  assign t[70] = (~t[95] & t[96]);
  assign t[71] = (~t[97] & t[98]);
  assign t[72] = (~t[99] & t[100]);
  assign t[73] = t[101] ^ x[2];
  assign t[74] = t[102] ^ x[3];
  assign t[75] = t[103] ^ x[5];
  assign t[76] = t[104] ^ x[6];
  assign t[77] = t[105] ^ x[8];
  assign t[78] = t[106] ^ x[9];
  assign t[79] = t[107] ^ x[11];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[108] ^ x[12];
  assign t[81] = t[109] ^ x[14];
  assign t[82] = t[110] ^ x[15];
  assign t[83] = t[111] ^ x[17];
  assign t[84] = t[112] ^ x[18];
  assign t[85] = t[113] ^ x[20];
  assign t[86] = t[114] ^ x[21];
  assign t[87] = t[115] ^ x[23];
  assign t[88] = t[116] ^ x[24];
  assign t[89] = t[117] ^ x[26];
  assign t[8] = ~(x[0]);
  assign t[90] = t[118] ^ x[27];
  assign t[91] = t[119] ^ x[29];
  assign t[92] = t[120] ^ x[30];
  assign t[93] = t[121] ^ x[32];
  assign t[94] = t[122] ^ x[33];
  assign t[95] = t[123] ^ x[35];
  assign t[96] = t[124] ^ x[36];
  assign t[97] = t[125] ^ x[38];
  assign t[98] = t[126] ^ x[39];
  assign t[99] = t[127] ^ x[41];
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [42:0] x;
 output y;

 wire [128:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[128] ^ x[42];
  assign t[101] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[1]);
  assign t[103] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[4]);
  assign t[105] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[7]);
  assign t[107] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[10]);
  assign t[109] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[13]);
  assign t[111] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[16]);
  assign t[113] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[19]);
  assign t[115] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[22]);
  assign t[117] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[25]);
  assign t[119] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[31]);
  assign t[120] = (x[28]);
  assign t[121] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[31]);
  assign t[123] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[34]);
  assign t[125] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[37]);
  assign t[127] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[40]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[32] | t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[33] & t[34]);
  assign t[16] = ~(t[35] & t[36]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[37] & t[8]);
  assign t[19] = ~(t[38] & t[39]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[40] & t[41]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[26] | t[31]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[26] & t[29]);
  assign t[26] = ~(t[44]);
  assign t[27] = ~(t[26] & t[30]);
  assign t[28] = ~(t[42] & t[11]);
  assign t[29] = t[22] & t[31];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[43]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = t[59] ^ x[3];
  assign t[46] = t[60] ^ x[6];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[15];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[21];
  assign t[52] = t[66] ^ x[24];
  assign t[53] = t[67] ^ x[27];
  assign t[54] = t[68] ^ x[30];
  assign t[55] = t[69] ^ x[33];
  assign t[56] = t[70] ^ x[36];
  assign t[57] = t[71] ^ x[39];
  assign t[58] = t[72] ^ x[42];
  assign t[59] = (~t[73] & t[74]);
  assign t[5] = ~(t[11]);
  assign t[60] = (~t[75] & t[76]);
  assign t[61] = (~t[77] & t[78]);
  assign t[62] = (~t[79] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[87] & t[88]);
  assign t[67] = (~t[89] & t[90]);
  assign t[68] = (~t[91] & t[92]);
  assign t[69] = (~t[93] & t[94]);
  assign t[6] = ~(t[12]);
  assign t[70] = (~t[95] & t[96]);
  assign t[71] = (~t[97] & t[98]);
  assign t[72] = (~t[99] & t[100]);
  assign t[73] = t[101] ^ x[2];
  assign t[74] = t[102] ^ x[3];
  assign t[75] = t[103] ^ x[5];
  assign t[76] = t[104] ^ x[6];
  assign t[77] = t[105] ^ x[8];
  assign t[78] = t[106] ^ x[9];
  assign t[79] = t[107] ^ x[11];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[108] ^ x[12];
  assign t[81] = t[109] ^ x[14];
  assign t[82] = t[110] ^ x[15];
  assign t[83] = t[111] ^ x[17];
  assign t[84] = t[112] ^ x[18];
  assign t[85] = t[113] ^ x[20];
  assign t[86] = t[114] ^ x[21];
  assign t[87] = t[115] ^ x[23];
  assign t[88] = t[116] ^ x[24];
  assign t[89] = t[117] ^ x[26];
  assign t[8] = ~(x[0]);
  assign t[90] = t[118] ^ x[27];
  assign t[91] = t[119] ^ x[29];
  assign t[92] = t[120] ^ x[30];
  assign t[93] = t[121] ^ x[32];
  assign t[94] = t[122] ^ x[33];
  assign t[95] = t[123] ^ x[35];
  assign t[96] = t[124] ^ x[36];
  assign t[97] = t[125] ^ x[38];
  assign t[98] = t[126] ^ x[39];
  assign t[99] = t[127] ^ x[41];
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[22]);
  assign t[103] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[25]);
  assign t[105] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[28]);
  assign t[107] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[31]);
  assign t[109] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[63] & t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (~t[65] & t[66]);
  assign t[51] = (~t[67] & t[68]);
  assign t[52] = (~t[69] & t[70]);
  assign t[53] = (~t[71] & t[72]);
  assign t[54] = (~t[73] & t[74]);
  assign t[55] = (~t[75] & t[76]);
  assign t[56] = (~t[77] & t[78]);
  assign t[57] = (~t[79] & t[80]);
  assign t[58] = (~t[81] & t[82]);
  assign t[59] = (~t[83] & t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (~t[85] & t[86]);
  assign t[61] = t[87] ^ x[1];
  assign t[62] = t[88] ^ x[2];
  assign t[63] = t[89] ^ x[5];
  assign t[64] = t[90] ^ x[6];
  assign t[65] = t[91] ^ x[8];
  assign t[66] = t[92] ^ x[9];
  assign t[67] = t[93] ^ x[11];
  assign t[68] = t[94] ^ x[12];
  assign t[69] = t[95] ^ x[14];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[15];
  assign t[71] = t[97] ^ x[17];
  assign t[72] = t[98] ^ x[18];
  assign t[73] = t[99] ^ x[20];
  assign t[74] = t[100] ^ x[21];
  assign t[75] = t[101] ^ x[23];
  assign t[76] = t[102] ^ x[24];
  assign t[77] = t[103] ^ x[26];
  assign t[78] = t[104] ^ x[27];
  assign t[79] = t[105] ^ x[29];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[30];
  assign t[81] = t[107] ^ x[32];
  assign t[82] = t[108] ^ x[33];
  assign t[83] = t[109] ^ x[35];
  assign t[84] = t[110] ^ x[36];
  assign t[85] = t[111] ^ x[38];
  assign t[86] = t[112] ^ x[39];
  assign t[87] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[0]);
  assign t[89] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[7]);
  assign t[93] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[10]);
  assign t[95] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[13]);
  assign t[97] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[16]);
  assign t[99] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind31(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind34(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[22]);
  assign t[103] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[25]);
  assign t[105] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[28]);
  assign t[107] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[31]);
  assign t[109] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[63] & t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (~t[65] & t[66]);
  assign t[51] = (~t[67] & t[68]);
  assign t[52] = (~t[69] & t[70]);
  assign t[53] = (~t[71] & t[72]);
  assign t[54] = (~t[73] & t[74]);
  assign t[55] = (~t[75] & t[76]);
  assign t[56] = (~t[77] & t[78]);
  assign t[57] = (~t[79] & t[80]);
  assign t[58] = (~t[81] & t[82]);
  assign t[59] = (~t[83] & t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (~t[85] & t[86]);
  assign t[61] = t[87] ^ x[1];
  assign t[62] = t[88] ^ x[2];
  assign t[63] = t[89] ^ x[5];
  assign t[64] = t[90] ^ x[6];
  assign t[65] = t[91] ^ x[8];
  assign t[66] = t[92] ^ x[9];
  assign t[67] = t[93] ^ x[11];
  assign t[68] = t[94] ^ x[12];
  assign t[69] = t[95] ^ x[14];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[15];
  assign t[71] = t[97] ^ x[17];
  assign t[72] = t[98] ^ x[18];
  assign t[73] = t[99] ^ x[20];
  assign t[74] = t[100] ^ x[21];
  assign t[75] = t[101] ^ x[23];
  assign t[76] = t[102] ^ x[24];
  assign t[77] = t[103] ^ x[26];
  assign t[78] = t[104] ^ x[27];
  assign t[79] = t[105] ^ x[29];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[30];
  assign t[81] = t[107] ^ x[32];
  assign t[82] = t[108] ^ x[33];
  assign t[83] = t[109] ^ x[35];
  assign t[84] = t[110] ^ x[36];
  assign t[85] = t[111] ^ x[38];
  assign t[86] = t[112] ^ x[39];
  assign t[87] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[0]);
  assign t[89] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[7]);
  assign t[93] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[10]);
  assign t[95] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[13]);
  assign t[97] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[16]);
  assign t[99] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[60] & t[61]);
  assign t[44] = (~t[62] & t[63]);
  assign t[45] = (~t[64] & t[65]);
  assign t[46] = (~t[66] & t[67]);
  assign t[47] = (~t[68] & t[69]);
  assign t[48] = t[70] ^ x[1];
  assign t[49] = t[71] ^ x[2];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[4];
  assign t[51] = t[73] ^ x[5];
  assign t[52] = t[74] ^ x[8];
  assign t[53] = t[75] ^ x[9];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[12];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[15];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[18];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[21];
  assign t[62] = t[84] ^ x[23];
  assign t[63] = t[85] ^ x[24];
  assign t[64] = t[86] ^ x[26];
  assign t[65] = t[87] ^ x[27];
  assign t[66] = t[88] ^ x[29];
  assign t[67] = t[89] ^ x[30];
  assign t[68] = t[90] ^ x[32];
  assign t[69] = t[91] ^ x[33];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[0]);
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[7]);
  assign t[76] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[10]);
  assign t[78] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[16]);
  assign t[82] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[19]);
  assign t[84] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[22]);
  assign t[86] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[25]);
  assign t[88] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind36(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind37(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind38(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind39(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[60] & t[61]);
  assign t[44] = (~t[62] & t[63]);
  assign t[45] = (~t[64] & t[65]);
  assign t[46] = (~t[66] & t[67]);
  assign t[47] = (~t[68] & t[69]);
  assign t[48] = t[70] ^ x[1];
  assign t[49] = t[71] ^ x[2];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[4];
  assign t[51] = t[73] ^ x[5];
  assign t[52] = t[74] ^ x[8];
  assign t[53] = t[75] ^ x[9];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[12];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[15];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[18];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[21];
  assign t[62] = t[84] ^ x[23];
  assign t[63] = t[85] ^ x[24];
  assign t[64] = t[86] ^ x[26];
  assign t[65] = t[87] ^ x[27];
  assign t[66] = t[88] ^ x[29];
  assign t[67] = t[89] ^ x[30];
  assign t[68] = t[90] ^ x[32];
  assign t[69] = t[91] ^ x[33];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[0]);
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[7]);
  assign t[76] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[10]);
  assign t[78] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[16]);
  assign t[82] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[19]);
  assign t[84] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[22]);
  assign t[86] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[25]);
  assign t[88] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = (~t[60] & t[61]);
  assign t[43] = (~t[62] & t[63]);
  assign t[44] = t[64] ^ x[1];
  assign t[45] = t[65] ^ x[2];
  assign t[46] = t[66] ^ x[4];
  assign t[47] = t[67] ^ x[5];
  assign t[48] = t[68] ^ x[8];
  assign t[49] = t[69] ^ x[9];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[11];
  assign t[51] = t[71] ^ x[12];
  assign t[52] = t[72] ^ x[14];
  assign t[53] = t[73] ^ x[15];
  assign t[54] = t[74] ^ x[17];
  assign t[55] = t[75] ^ x[18];
  assign t[56] = t[76] ^ x[20];
  assign t[57] = t[77] ^ x[21];
  assign t[58] = t[78] ^ x[23];
  assign t[59] = t[79] ^ x[24];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[26];
  assign t[61] = t[81] ^ x[27];
  assign t[62] = t[82] ^ x[29];
  assign t[63] = t[83] ^ x[30];
  assign t[64] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[0]);
  assign t[66] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[3]);
  assign t[68] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[10]);
  assign t[72] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[13]);
  assign t[74] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[16]);
  assign t[76] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[19]);
  assign t[78] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[25]);
  assign t[82] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind41(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind42(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind43(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind44(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = (~t[60] & t[61]);
  assign t[43] = (~t[62] & t[63]);
  assign t[44] = t[64] ^ x[1];
  assign t[45] = t[65] ^ x[2];
  assign t[46] = t[66] ^ x[4];
  assign t[47] = t[67] ^ x[5];
  assign t[48] = t[68] ^ x[8];
  assign t[49] = t[69] ^ x[9];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[11];
  assign t[51] = t[71] ^ x[12];
  assign t[52] = t[72] ^ x[14];
  assign t[53] = t[73] ^ x[15];
  assign t[54] = t[74] ^ x[17];
  assign t[55] = t[75] ^ x[18];
  assign t[56] = t[76] ^ x[20];
  assign t[57] = t[77] ^ x[21];
  assign t[58] = t[78] ^ x[23];
  assign t[59] = t[79] ^ x[24];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[26];
  assign t[61] = t[81] ^ x[27];
  assign t[62] = t[82] ^ x[29];
  assign t[63] = t[83] ^ x[30];
  assign t[64] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[0]);
  assign t[66] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[3]);
  assign t[68] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[10]);
  assign t[72] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[13]);
  assign t[74] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[16]);
  assign t[76] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[19]);
  assign t[78] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[25]);
  assign t[82] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = (~t[54] & t[55]);
  assign t[39] = (~t[56] & t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[1];
  assign t[41] = t[59] ^ x[2];
  assign t[42] = t[60] ^ x[5];
  assign t[43] = t[61] ^ x[6];
  assign t[44] = t[62] ^ x[8];
  assign t[45] = t[63] ^ x[9];
  assign t[46] = t[64] ^ x[11];
  assign t[47] = t[65] ^ x[12];
  assign t[48] = t[66] ^ x[14];
  assign t[49] = t[67] ^ x[15];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[17];
  assign t[51] = t[69] ^ x[18];
  assign t[52] = t[70] ^ x[20];
  assign t[53] = t[71] ^ x[21];
  assign t[54] = t[72] ^ x[23];
  assign t[55] = t[73] ^ x[24];
  assign t[56] = t[74] ^ x[26];
  assign t[57] = t[75] ^ x[27];
  assign t[58] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[4]);
  assign t[62] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[7]);
  assign t[64] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[10]);
  assign t[66] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[13]);
  assign t[68] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[19]);
  assign t[72] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[22]);
  assign t[74] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind46(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind47(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind48(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind49(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = (~t[54] & t[55]);
  assign t[39] = (~t[56] & t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[1];
  assign t[41] = t[59] ^ x[2];
  assign t[42] = t[60] ^ x[5];
  assign t[43] = t[61] ^ x[6];
  assign t[44] = t[62] ^ x[8];
  assign t[45] = t[63] ^ x[9];
  assign t[46] = t[64] ^ x[11];
  assign t[47] = t[65] ^ x[12];
  assign t[48] = t[66] ^ x[14];
  assign t[49] = t[67] ^ x[15];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[17];
  assign t[51] = t[69] ^ x[18];
  assign t[52] = t[70] ^ x[20];
  assign t[53] = t[71] ^ x[21];
  assign t[54] = t[72] ^ x[23];
  assign t[55] = t[73] ^ x[24];
  assign t[56] = t[74] ^ x[26];
  assign t[57] = t[75] ^ x[27];
  assign t[58] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[4]);
  assign t[62] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[7]);
  assign t[64] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[10]);
  assign t[66] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[13]);
  assign t[68] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[19]);
  assign t[72] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[22]);
  assign t[74] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = (~t[73] & t[74]);
  assign t[52] = (~t[75] & t[76]);
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[6];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[9];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[12];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[15];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[18];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[21];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[24];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[27];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[30];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[33];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[36];
  assign t[77] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[0]);
  assign t[79] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[7]);
  assign t[83] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[10]);
  assign t[85] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[13]);
  assign t[87] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[16]);
  assign t[89] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[22]);
  assign t[93] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[25]);
  assign t[95] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[28]);
  assign t[97] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[31]);
  assign t[99] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind51(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind52(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind53(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind54(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = (~t[73] & t[74]);
  assign t[52] = (~t[75] & t[76]);
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[6];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[9];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[12];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[15];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[18];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[21];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[24];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[27];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[30];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[33];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[36];
  assign t[77] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[0]);
  assign t[79] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[7]);
  assign t[83] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[10]);
  assign t[85] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[13]);
  assign t[87] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[16]);
  assign t[89] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[22]);
  assign t[93] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[25]);
  assign t[95] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[28]);
  assign t[97] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[31]);
  assign t[99] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[20]);
  assign t[13] = t[14] & t[21];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = t[15] ^ t[4];
  assign t[30] = t[39] ^ x[20];
  assign t[31] = t[40] ^ x[23];
  assign t[32] = t[41] ^ x[26];
  assign t[33] = (~t[42] & t[43]);
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = ~(t[16]);
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = t[60] ^ x[1];
  assign t[43] = t[61] ^ x[2];
  assign t[44] = t[62] ^ x[4];
  assign t[45] = t[63] ^ x[5];
  assign t[46] = t[64] ^ x[7];
  assign t[47] = t[65] ^ x[8];
  assign t[48] = t[66] ^ x[10];
  assign t[49] = t[67] ^ x[11];
  assign t[4] = ~(t[5] & t[17]);
  assign t[50] = t[68] ^ x[13];
  assign t[51] = t[69] ^ x[14];
  assign t[52] = t[70] ^ x[16];
  assign t[53] = t[71] ^ x[17];
  assign t[54] = t[72] ^ x[19];
  assign t[55] = t[73] ^ x[20];
  assign t[56] = t[74] ^ x[22];
  assign t[57] = t[75] ^ x[23];
  assign t[58] = t[76] ^ x[25];
  assign t[59] = t[77] ^ x[26];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[0]);
  assign t[62] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[3]);
  assign t[64] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[6]);
  assign t[66] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[9]);
  assign t[68] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[12]);
  assign t[6] = ~(t[18]);
  assign t[70] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[15]);
  assign t[72] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[18]);
  assign t[74] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[21]);
  assign t[76] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[19] | t[10]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind56(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind57(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind58(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind59(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[20]);
  assign t[13] = t[14] & t[21];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = t[15] ^ t[4];
  assign t[30] = t[39] ^ x[20];
  assign t[31] = t[40] ^ x[23];
  assign t[32] = t[41] ^ x[26];
  assign t[33] = (~t[42] & t[43]);
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = ~(t[16]);
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = t[60] ^ x[1];
  assign t[43] = t[61] ^ x[2];
  assign t[44] = t[62] ^ x[4];
  assign t[45] = t[63] ^ x[5];
  assign t[46] = t[64] ^ x[7];
  assign t[47] = t[65] ^ x[8];
  assign t[48] = t[66] ^ x[10];
  assign t[49] = t[67] ^ x[11];
  assign t[4] = ~(t[5] & t[17]);
  assign t[50] = t[68] ^ x[13];
  assign t[51] = t[69] ^ x[14];
  assign t[52] = t[70] ^ x[16];
  assign t[53] = t[71] ^ x[17];
  assign t[54] = t[72] ^ x[19];
  assign t[55] = t[73] ^ x[20];
  assign t[56] = t[74] ^ x[22];
  assign t[57] = t[75] ^ x[23];
  assign t[58] = t[76] ^ x[25];
  assign t[59] = t[77] ^ x[26];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[0]);
  assign t[62] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[3]);
  assign t[64] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[6]);
  assign t[66] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[9]);
  assign t[68] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[12]);
  assign t[6] = ~(t[18]);
  assign t[70] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[15]);
  assign t[72] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[18]);
  assign t[74] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[21]);
  assign t[76] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[19] | t[10]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [29:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[22] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[23]);
  assign t[15] = t[16] & t[24];
  assign t[16] = ~(t[25] | t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[17] ^ t[3]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = t[37] ^ x[2];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = (~t[47] & t[48]);
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = t[67] ^ x[1];
  assign t[48] = t[68] ^ x[2];
  assign t[49] = t[69] ^ x[4];
  assign t[4] = ~(t[18]);
  assign t[50] = t[70] ^ x[5];
  assign t[51] = t[71] ^ x[7];
  assign t[52] = t[72] ^ x[8];
  assign t[53] = t[73] ^ x[10];
  assign t[54] = t[74] ^ x[11];
  assign t[55] = t[75] ^ x[13];
  assign t[56] = t[76] ^ x[14];
  assign t[57] = t[77] ^ x[16];
  assign t[58] = t[78] ^ x[17];
  assign t[59] = t[79] ^ x[19];
  assign t[5] = ~(t[19]);
  assign t[60] = t[80] ^ x[20];
  assign t[61] = t[81] ^ x[22];
  assign t[62] = t[82] ^ x[23];
  assign t[63] = t[83] ^ x[25];
  assign t[64] = t[84] ^ x[26];
  assign t[65] = t[85] ^ x[28];
  assign t[66] = t[86] ^ x[29];
  assign t[67] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[0]);
  assign t[69] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[7] & t[20]);
  assign t[70] = (x[3]);
  assign t[71] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[6]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[8] | t[9]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[21]);
  assign t[83] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[24]);
  assign t[85] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[27]);
  assign t[8] = ~(t[21]);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind61(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind62(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind63(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind64(x, y);
 input [29:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[22] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[23]);
  assign t[15] = t[16] & t[24];
  assign t[16] = ~(t[25] | t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[17] ^ t[3]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = t[37] ^ x[2];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = (~t[47] & t[48]);
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = t[67] ^ x[1];
  assign t[48] = t[68] ^ x[2];
  assign t[49] = t[69] ^ x[4];
  assign t[4] = ~(t[18]);
  assign t[50] = t[70] ^ x[5];
  assign t[51] = t[71] ^ x[7];
  assign t[52] = t[72] ^ x[8];
  assign t[53] = t[73] ^ x[10];
  assign t[54] = t[74] ^ x[11];
  assign t[55] = t[75] ^ x[13];
  assign t[56] = t[76] ^ x[14];
  assign t[57] = t[77] ^ x[16];
  assign t[58] = t[78] ^ x[17];
  assign t[59] = t[79] ^ x[19];
  assign t[5] = ~(t[19]);
  assign t[60] = t[80] ^ x[20];
  assign t[61] = t[81] ^ x[22];
  assign t[62] = t[82] ^ x[23];
  assign t[63] = t[83] ^ x[25];
  assign t[64] = t[84] ^ x[26];
  assign t[65] = t[85] ^ x[28];
  assign t[66] = t[86] ^ x[29];
  assign t[67] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[0]);
  assign t[69] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[7] & t[20]);
  assign t[70] = (x[3]);
  assign t[71] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[6]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[8] | t[9]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[21]);
  assign t[83] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[24]);
  assign t[85] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[27]);
  assign t[8] = ~(t[21]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[18]);
  assign t[12] = t[13] & t[19];
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[4]);
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[2];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[5];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[8];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[11];
  assign t[46] = t[62] ^ x[13];
  assign t[47] = t[63] ^ x[14];
  assign t[48] = t[64] ^ x[16];
  assign t[49] = t[65] ^ x[17];
  assign t[4] = ~(t[15]);
  assign t[50] = t[66] ^ x[19];
  assign t[51] = t[67] ^ x[20];
  assign t[52] = t[68] ^ x[22];
  assign t[53] = t[69] ^ x[23];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[16]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[17] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind66(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind67(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind68(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind69(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[18]);
  assign t[12] = t[13] & t[19];
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[4]);
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[2];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[5];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[8];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[11];
  assign t[46] = t[62] ^ x[13];
  assign t[47] = t[63] ^ x[14];
  assign t[48] = t[64] ^ x[16];
  assign t[49] = t[65] ^ x[17];
  assign t[4] = ~(t[15]);
  assign t[50] = t[66] ^ x[19];
  assign t[51] = t[67] ^ x[20];
  assign t[52] = t[68] ^ x[22];
  assign t[53] = t[69] ^ x[23];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[16]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[17] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [20:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[11] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = t[26] ^ x[2];
  assign t[1] = ~(t[3]);
  assign t[20] = t[27] ^ x[5];
  assign t[21] = t[28] ^ x[8];
  assign t[22] = t[29] ^ x[11];
  assign t[23] = t[30] ^ x[14];
  assign t[24] = t[31] ^ x[17];
  assign t[25] = t[32] ^ x[20];
  assign t[26] = (~t[33] & t[34]);
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = t[47] ^ x[1];
  assign t[34] = t[48] ^ x[2];
  assign t[35] = t[49] ^ x[4];
  assign t[36] = t[50] ^ x[5];
  assign t[37] = t[51] ^ x[7];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[10];
  assign t[3] = ~(t[12]);
  assign t[40] = t[54] ^ x[11];
  assign t[41] = t[55] ^ x[13];
  assign t[42] = t[56] ^ x[14];
  assign t[43] = t[57] ^ x[16];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[19];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[48] = (x[0]);
  assign t[49] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[13]);
  assign t[50] = (x[3]);
  assign t[51] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[6]);
  assign t[53] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[9]);
  assign t[55] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[12]);
  assign t[57] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[15]);
  assign t[59] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[18]);
  assign t[6] = ~(t[14] | t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind71(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind72(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind73(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind74(x, y);
 input [20:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[11] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = t[26] ^ x[2];
  assign t[1] = ~(t[3]);
  assign t[20] = t[27] ^ x[5];
  assign t[21] = t[28] ^ x[8];
  assign t[22] = t[29] ^ x[11];
  assign t[23] = t[30] ^ x[14];
  assign t[24] = t[31] ^ x[17];
  assign t[25] = t[32] ^ x[20];
  assign t[26] = (~t[33] & t[34]);
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = t[47] ^ x[1];
  assign t[34] = t[48] ^ x[2];
  assign t[35] = t[49] ^ x[4];
  assign t[36] = t[50] ^ x[5];
  assign t[37] = t[51] ^ x[7];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[10];
  assign t[3] = ~(t[12]);
  assign t[40] = t[54] ^ x[11];
  assign t[41] = t[55] ^ x[13];
  assign t[42] = t[56] ^ x[14];
  assign t[43] = t[57] ^ x[16];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[19];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[48] = (x[0]);
  assign t[49] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[13]);
  assign t[50] = (x[3]);
  assign t[51] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[6]);
  assign t[53] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[9]);
  assign t[55] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[12]);
  assign t[57] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[15]);
  assign t[59] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[18]);
  assign t[6] = ~(t[14] | t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [11:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[5] | t[1]);
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (~t[17] & t[18]);
  assign t[14] = (~t[19] & t[20]);
  assign t[15] = (~t[21] & t[22]);
  assign t[16] = (~t[23] & t[24]);
  assign t[17] = t[25] ^ x[1];
  assign t[18] = t[26] ^ x[2];
  assign t[19] = t[27] ^ x[4];
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[7];
  assign t[22] = t[30] ^ x[8];
  assign t[23] = t[31] ^ x[10];
  assign t[24] = t[32] ^ x[11];
  assign t[25] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[0]);
  assign t[27] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[3]);
  assign t[29] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (x[6]);
  assign t[31] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~(t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind76(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind77(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind78(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind79(x, y);
 input [11:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[5] | t[1]);
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (~t[17] & t[18]);
  assign t[14] = (~t[19] & t[20]);
  assign t[15] = (~t[21] & t[22]);
  assign t[16] = (~t[23] & t[24]);
  assign t[17] = t[25] ^ x[1];
  assign t[18] = t[26] ^ x[2];
  assign t[19] = t[27] ^ x[4];
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[7];
  assign t[22] = t[30] ^ x[8];
  assign t[23] = t[31] ^ x[10];
  assign t[24] = t[32] ^ x[11];
  assign t[25] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[0]);
  assign t[27] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[3]);
  assign t[29] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (x[6]);
  assign t[31] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~(t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [12:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[3];
  assign t[14] = t[18] ^ x[6];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[11];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(x[0]);
  assign t[30] = (x[1]);
  assign t[31] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[4]);
  assign t[33] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[7]);
  assign t[35] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind81(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind82(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind83(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind84(x, y);
 input [12:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[3];
  assign t[14] = t[18] ^ x[6];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[3];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[6];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[11];
  assign t[28] = t[36] ^ x[12];
  assign t[29] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(x[0]);
  assign t[30] = (x[1]);
  assign t[31] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[4]);
  assign t[33] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[7]);
  assign t[35] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = t[20] ^ x[2];
  assign t[15] = t[21] ^ x[5];
  assign t[16] = t[22] ^ x[8];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = ~(t[8] | t[3]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = (~t[34] & t[35]);
  assign t[25] = (~t[36] & t[37]);
  assign t[26] = t[38] ^ x[1];
  assign t[27] = t[39] ^ x[2];
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[9]);
  assign t[30] = t[42] ^ x[7];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[10];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[13];
  assign t[35] = t[47] ^ x[14];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[17];
  assign t[38] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[0]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[3]);
  assign t[42] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[6]);
  assign t[44] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[9]);
  assign t[46] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[12]);
  assign t[48] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[15]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = t[7] & t[11];
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind86(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind87(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind88(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind89(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = t[20] ^ x[2];
  assign t[15] = t[21] ^ x[5];
  assign t[16] = t[22] ^ x[8];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = ~(t[8] | t[3]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = (~t[34] & t[35]);
  assign t[25] = (~t[36] & t[37]);
  assign t[26] = t[38] ^ x[1];
  assign t[27] = t[39] ^ x[2];
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[9]);
  assign t[30] = t[42] ^ x[7];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[10];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[13];
  assign t[35] = t[47] ^ x[14];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[17];
  assign t[38] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[0]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[3]);
  assign t[42] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[6]);
  assign t[44] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[9]);
  assign t[46] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[12]);
  assign t[48] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[15]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = t[7] & t[11];
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind91(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind92(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind93(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind94(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind96(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind97(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind98(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind99(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind101(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind102(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind103(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind104(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind106(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind107(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind108(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind109(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind111(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind112(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind113(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind114(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind116(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind117(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind118(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind119(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind121(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind122(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind123(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind124(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind126(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind127(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind128(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind129(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind131(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind132(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind133(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind134(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[1];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [67:0] x;
 output y;

 wire [190:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[57];
  assign t[101] = t[123] ^ x[58];
  assign t[102] = t[124] ^ x[64];
  assign t[103] = t[125] ^ x[66];
  assign t[104] = t[126] ^ x[67];
  assign t[105] = (~t[127] & t[128]);
  assign t[106] = (~t[129] & t[130]);
  assign t[107] = (~t[131] & t[132]);
  assign t[108] = (~t[133] & t[134]);
  assign t[109] = (~t[135] & t[136]);
  assign t[10] = t[65] ^ t[66];
  assign t[110] = (~t[137] & t[138]);
  assign t[111] = (~t[139] & t[140]);
  assign t[112] = (~t[139] & t[141]);
  assign t[113] = (~t[139] & t[142]);
  assign t[114] = (~t[139] & t[143]);
  assign t[115] = (~t[129] & t[144]);
  assign t[116] = (~t[145] & t[146]);
  assign t[117] = (~t[135] & t[147]);
  assign t[118] = (~t[137] & t[148]);
  assign t[119] = (~t[129] & t[149]);
  assign t[11] = ~(t[14]);
  assign t[120] = (~t[150] & t[151]);
  assign t[121] = (~t[135] & t[152]);
  assign t[122] = (~t[137] & t[153]);
  assign t[123] = (~t[129] & t[154]);
  assign t[124] = (~t[155] & t[156]);
  assign t[125] = (~t[135] & t[157]);
  assign t[126] = (~t[137] & t[158]);
  assign t[127] = t[159] ^ x[1];
  assign t[128] = t[160] ^ x[2];
  assign t[129] = t[161] ^ x[7];
  assign t[12] = ~(t[15] | t[67]);
  assign t[130] = t[162] ^ x[8];
  assign t[131] = t[163] ^ x[10];
  assign t[132] = t[164] ^ x[11];
  assign t[133] = t[165] ^ x[13];
  assign t[134] = t[166] ^ x[14];
  assign t[135] = t[167] ^ x[20];
  assign t[136] = t[168] ^ x[21];
  assign t[137] = t[169] ^ x[26];
  assign t[138] = t[170] ^ x[27];
  assign t[139] = t[171] ^ x[32];
  assign t[13] = ~(t[68] ^ t[69]);
  assign t[140] = t[172] ^ x[33];
  assign t[141] = t[173] ^ x[34];
  assign t[142] = t[174] ^ x[35];
  assign t[143] = t[175] ^ x[37];
  assign t[144] = t[176] ^ x[38];
  assign t[145] = t[177] ^ x[43];
  assign t[146] = t[178] ^ x[44];
  assign t[147] = t[179] ^ x[46];
  assign t[148] = t[180] ^ x[47];
  assign t[149] = t[181] ^ x[48];
  assign t[14] = ~(x[36]);
  assign t[150] = t[182] ^ x[53];
  assign t[151] = t[183] ^ x[54];
  assign t[152] = t[184] ^ x[56];
  assign t[153] = t[185] ^ x[57];
  assign t[154] = t[186] ^ x[58];
  assign t[155] = t[187] ^ x[63];
  assign t[156] = t[188] ^ x[64];
  assign t[157] = t[189] ^ x[66];
  assign t[158] = t[190] ^ x[67];
  assign t[159] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = ~(t[70]);
  assign t[160] = (x[0]);
  assign t[161] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[162] = (x[3]);
  assign t[163] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[164] = (x[9]);
  assign t[165] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[166] = (x[12]);
  assign t[167] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[16] = ~(t[17] & t[18]);
  assign t[170] = (x[25]);
  assign t[171] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[172] = (x[29]);
  assign t[173] = (x[31]);
  assign t[174] = (x[28]);
  assign t[175] = (x[30]);
  assign t[176] = (x[4]);
  assign t[177] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[18]);
  assign t[17] = t[61] ? t[20] : t[19];
  assign t[180] = (x[24]);
  assign t[181] = (x[5]);
  assign t[182] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[17]);
  assign t[185] = (x[23]);
  assign t[186] = (x[6]);
  assign t[187] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[188] = (x[62]);
  assign t[189] = (x[16]);
  assign t[18] = ~(t[5] & t[21]);
  assign t[190] = (x[22]);
  assign t[19] = ~(t[71]);
  assign t[1] = t[61] ? t[4] : t[3];
  assign t[20] = ~(t[63] & t[22]);
  assign t[21] = t[64] ? t[24] : t[23];
  assign t[22] = t[11] ? x[45] : t[72];
  assign t[23] = ~(t[25] | t[26]);
  assign t[24] = t[73] ^ t[74];
  assign t[25] = ~(t[27] | t[28]);
  assign t[26] = ~(t[15] | t[13]);
  assign t[27] = ~(t[29] | t[15]);
  assign t[28] = t[68] ? t[30] : t[67];
  assign t[29] = ~(t[68] | t[69]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[67] & t[31]);
  assign t[31] = ~(t[32] & t[15]);
  assign t[32] = ~(t[69]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[61] ? t[37] : t[36];
  assign t[35] = ~(t[5] & t[38]);
  assign t[36] = ~(t[75]);
  assign t[37] = ~(t[63] & t[39]);
  assign t[38] = t[64] ? t[41] : t[40];
  assign t[39] = t[11] ? x[55] : t[76];
  assign t[3] = ~(t[62]);
  assign t[40] = ~(t[42] & t[43]);
  assign t[41] = t[77] ^ t[78];
  assign t[42] = ~(t[44] & t[30]);
  assign t[43] = ~(t[27] & t[28]);
  assign t[44] = ~(t[70] | t[45]);
  assign t[45] = ~(t[46] | t[47]);
  assign t[46] = ~(t[68]);
  assign t[47] = ~(t[32] & t[48]);
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[50] & t[51]);
  assign t[4] = ~(t[63] & t[7]);
  assign t[50] = t[61] ? t[53] : t[52];
  assign t[51] = ~(t[5] & t[54]);
  assign t[52] = ~(t[79]);
  assign t[53] = ~(t[63] & t[55]);
  assign t[54] = t[64] ? t[57] : t[56];
  assign t[55] = t[11] ? x[65] : t[80];
  assign t[56] = ~(t[58] & t[59]);
  assign t[57] = t[81] ^ t[82];
  assign t[58] = t[68] ? t[60] : t[30];
  assign t[59] = ~(t[29] & t[48]);
  assign t[5] = ~(t[63] | t[8]);
  assign t[60] = ~(t[15] & t[47]);
  assign t[61] = (t[83]);
  assign t[62] = (t[84]);
  assign t[63] = (t[85]);
  assign t[64] = (t[86]);
  assign t[65] = (t[87]);
  assign t[66] = (t[88]);
  assign t[67] = (t[89]);
  assign t[68] = (t[90]);
  assign t[69] = (t[91]);
  assign t[6] = t[64] ? t[10] : t[9];
  assign t[70] = (t[92]);
  assign t[71] = (t[93]);
  assign t[72] = (t[94]);
  assign t[73] = (t[95]);
  assign t[74] = (t[96]);
  assign t[75] = (t[97]);
  assign t[76] = (t[98]);
  assign t[77] = (t[99]);
  assign t[78] = (t[100]);
  assign t[79] = (t[101]);
  assign t[7] = t[11] ? x[15] : t[62];
  assign t[80] = (t[102]);
  assign t[81] = (t[103]);
  assign t[82] = (t[104]);
  assign t[83] = t[105] ^ x[2];
  assign t[84] = t[106] ^ x[8];
  assign t[85] = t[107] ^ x[11];
  assign t[86] = t[108] ^ x[14];
  assign t[87] = t[109] ^ x[21];
  assign t[88] = t[110] ^ x[27];
  assign t[89] = t[111] ^ x[33];
  assign t[8] = ~(t[61]);
  assign t[90] = t[112] ^ x[34];
  assign t[91] = t[113] ^ x[35];
  assign t[92] = t[114] ^ x[37];
  assign t[93] = t[115] ^ x[38];
  assign t[94] = t[116] ^ x[44];
  assign t[95] = t[117] ^ x[46];
  assign t[96] = t[118] ^ x[47];
  assign t[97] = t[119] ^ x[48];
  assign t[98] = t[120] ^ x[54];
  assign t[99] = t[121] ^ x[56];
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0] & ~t[16] & ~t[33] & ~t[49]) | (~t[0] & t[16] & ~t[33] & ~t[49]) | (~t[0] & ~t[16] & t[33] & ~t[49]) | (~t[0] & ~t[16] & ~t[33] & t[49]) | (t[0] & t[16] & t[33] & ~t[49]) | (t[0] & t[16] & ~t[33] & t[49]) | (t[0] & ~t[16] & t[33] & t[49]) | (~t[0] & t[16] & t[33] & t[49]);
endmodule

module R2ind136(x, y);
 input [43:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = t[30] ? t[16] : t[15];
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[40]);
  assign t[15] = ~(t[31] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[30] | t[32]);
  assign t[18] = ~(t[31]);
  assign t[19] = ~(t[22] & t[20]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[22] & t[18]);
  assign t[22] = ~(t[32]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[8];
  assign t[36] = t[47] ^ x[11];
  assign t[37] = t[48] ^ x[14];
  assign t[38] = t[49] ^ x[20];
  assign t[39] = t[50] ^ x[27];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[33];
  assign t[41] = t[52] ^ x[39];
  assign t[42] = t[53] ^ x[41];
  assign t[43] = t[54] ^ x[42];
  assign t[44] = t[55] ^ x[43];
  assign t[45] = (~t[56] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[60] & t[61]);
  assign t[48] = (~t[62] & t[63]);
  assign t[49] = (~t[64] & t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (~t[66] & t[67]);
  assign t[51] = (~t[68] & t[69]);
  assign t[52] = (~t[70] & t[71]);
  assign t[53] = (~t[70] & t[72]);
  assign t[54] = (~t[70] & t[73]);
  assign t[55] = (~t[70] & t[74]);
  assign t[56] = t[75] ^ x[1];
  assign t[57] = t[76] ^ x[2];
  assign t[58] = t[77] ^ x[7];
  assign t[59] = t[78] ^ x[8];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[79] ^ x[10];
  assign t[61] = t[80] ^ x[11];
  assign t[62] = t[81] ^ x[13];
  assign t[63] = t[82] ^ x[14];
  assign t[64] = t[83] ^ x[19];
  assign t[65] = t[84] ^ x[20];
  assign t[66] = t[85] ^ x[26];
  assign t[67] = t[86] ^ x[27];
  assign t[68] = t[87] ^ x[32];
  assign t[69] = t[88] ^ x[33];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[89] ^ x[38];
  assign t[71] = t[90] ^ x[39];
  assign t[72] = t[91] ^ x[41];
  assign t[73] = t[92] ^ x[42];
  assign t[74] = t[93] ^ x[43];
  assign t[75] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[0]);
  assign t[77] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[78] = (x[6]);
  assign t[79] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[11] ? x[21] : t[27];
  assign t[80] = (x[9]);
  assign t[81] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[12]);
  assign t[83] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[84] = (x[18]);
  assign t[85] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[86] = (x[22]);
  assign t[87] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[88] = (x[28]);
  assign t[89] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[37]);
  assign t[91] = (x[35]);
  assign t[92] = (x[34]);
  assign t[93] = (x[36]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [43:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[32] ^ t[33];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[34]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[35] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = t[36] ? t[16] : t[35];
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = t[27] ? t[4] : t[3];
  assign t[20] = ~(t[25] & t[22]);
  assign t[21] = ~(t[36] | t[37]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[36]);
  assign t[24] = ~(t[25] & t[26]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[35]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = (t[47]);
  assign t[37] = (t[48]);
  assign t[38] = t[49] ^ x[2];
  assign t[39] = t[50] ^ x[8];
  assign t[3] = ~(t[28]);
  assign t[40] = t[51] ^ x[11];
  assign t[41] = t[52] ^ x[14];
  assign t[42] = t[53] ^ x[20];
  assign t[43] = t[54] ^ x[27];
  assign t[44] = t[55] ^ x[33];
  assign t[45] = t[56] ^ x[40];
  assign t[46] = t[57] ^ x[41];
  assign t[47] = t[58] ^ x[42];
  assign t[48] = t[59] ^ x[43];
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[29] & t[7]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = (~t[66] & t[67]);
  assign t[53] = (~t[68] & t[69]);
  assign t[54] = (~t[70] & t[71]);
  assign t[55] = (~t[72] & t[73]);
  assign t[56] = (~t[74] & t[75]);
  assign t[57] = (~t[74] & t[76]);
  assign t[58] = (~t[74] & t[77]);
  assign t[59] = (~t[74] & t[78]);
  assign t[5] = ~(t[29] | t[8]);
  assign t[60] = t[79] ^ x[1];
  assign t[61] = t[80] ^ x[2];
  assign t[62] = t[81] ^ x[7];
  assign t[63] = t[82] ^ x[8];
  assign t[64] = t[83] ^ x[10];
  assign t[65] = t[84] ^ x[11];
  assign t[66] = t[85] ^ x[13];
  assign t[67] = t[86] ^ x[14];
  assign t[68] = t[87] ^ x[19];
  assign t[69] = t[88] ^ x[20];
  assign t[6] = t[30] ? t[10] : t[9];
  assign t[70] = t[89] ^ x[26];
  assign t[71] = t[90] ^ x[27];
  assign t[72] = t[91] ^ x[32];
  assign t[73] = t[92] ^ x[33];
  assign t[74] = t[93] ^ x[39];
  assign t[75] = t[94] ^ x[40];
  assign t[76] = t[95] ^ x[41];
  assign t[77] = t[96] ^ x[42];
  assign t[78] = t[97] ^ x[43];
  assign t[79] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[11] ? x[21] : t[31];
  assign t[80] = (x[0]);
  assign t[81] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[82] = (x[5]);
  assign t[83] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[9]);
  assign t[85] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[12]);
  assign t[87] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[88] = (x[18]);
  assign t[89] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[8] = ~(t[27]);
  assign t[90] = (x[23]);
  assign t[91] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[92] = (x[29]);
  assign t[93] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[94] = (x[37]);
  assign t[95] = (x[36]);
  assign t[96] = (x[38]);
  assign t[97] = (x[35]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [43:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(x[34]);
  assign t[15] = ~(t[19] | t[17]);
  assign t[16] = t[30] ? t[20] : t[31];
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[30] ^ t[33]);
  assign t[19] = ~(t[30] | t[33]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[31] & t[21]);
  assign t[21] = ~(t[22] & t[17]);
  assign t[22] = ~(t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[8];
  assign t[36] = t[47] ^ x[11];
  assign t[37] = t[48] ^ x[14];
  assign t[38] = t[49] ^ x[20];
  assign t[39] = t[50] ^ x[27];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[33];
  assign t[41] = t[52] ^ x[40];
  assign t[42] = t[53] ^ x[41];
  assign t[43] = t[54] ^ x[42];
  assign t[44] = t[55] ^ x[43];
  assign t[45] = (~t[56] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[60] & t[61]);
  assign t[48] = (~t[62] & t[63]);
  assign t[49] = (~t[64] & t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (~t[66] & t[67]);
  assign t[51] = (~t[68] & t[69]);
  assign t[52] = (~t[70] & t[71]);
  assign t[53] = (~t[70] & t[72]);
  assign t[54] = (~t[70] & t[73]);
  assign t[55] = (~t[70] & t[74]);
  assign t[56] = t[75] ^ x[1];
  assign t[57] = t[76] ^ x[2];
  assign t[58] = t[77] ^ x[7];
  assign t[59] = t[78] ^ x[8];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[79] ^ x[10];
  assign t[61] = t[80] ^ x[11];
  assign t[62] = t[81] ^ x[13];
  assign t[63] = t[82] ^ x[14];
  assign t[64] = t[83] ^ x[19];
  assign t[65] = t[84] ^ x[20];
  assign t[66] = t[85] ^ x[26];
  assign t[67] = t[86] ^ x[27];
  assign t[68] = t[87] ^ x[32];
  assign t[69] = t[88] ^ x[33];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[89] ^ x[39];
  assign t[71] = t[90] ^ x[40];
  assign t[72] = t[91] ^ x[41];
  assign t[73] = t[92] ^ x[42];
  assign t[74] = t[93] ^ x[43];
  assign t[75] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[0]);
  assign t[77] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[78] = (x[4]);
  assign t[79] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[11] ? x[21] : t[27];
  assign t[80] = (x[9]);
  assign t[81] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[12]);
  assign t[83] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[84] = (x[18]);
  assign t[85] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[86] = (x[24]);
  assign t[87] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[88] = (x[30]);
  assign t[89] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[38]);
  assign t[91] = (x[36]);
  assign t[92] = (x[37]);
  assign t[93] = (x[35]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [37:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[20] ^ t[21];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[22]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[14] = ~(x[36]);
  assign t[15] = ~(t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = t[16] ? t[4] : t[3];
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[11];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[27];
  assign t[32] = t[42] ^ x[33];
  assign t[33] = t[43] ^ x[34];
  assign t[34] = t[44] ^ x[35];
  assign t[35] = t[45] ^ x[37];
  assign t[36] = (~t[46] & t[47]);
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[17]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[58] & t[60]);
  assign t[44] = (~t[58] & t[61]);
  assign t[45] = (~t[58] & t[62]);
  assign t[46] = t[63] ^ x[1];
  assign t[47] = t[64] ^ x[2];
  assign t[48] = t[65] ^ x[7];
  assign t[49] = t[66] ^ x[8];
  assign t[4] = ~(t[18] & t[7]);
  assign t[50] = t[67] ^ x[10];
  assign t[51] = t[68] ^ x[11];
  assign t[52] = t[69] ^ x[13];
  assign t[53] = t[70] ^ x[14];
  assign t[54] = t[71] ^ x[20];
  assign t[55] = t[72] ^ x[21];
  assign t[56] = t[73] ^ x[26];
  assign t[57] = t[74] ^ x[27];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = ~(t[18] | t[8]);
  assign t[60] = t[77] ^ x[34];
  assign t[61] = t[78] ^ x[35];
  assign t[62] = t[79] ^ x[37];
  assign t[63] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[0]);
  assign t[65] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[66] = (x[3]);
  assign t[67] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[9]);
  assign t[69] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = t[19] ? t[10] : t[9];
  assign t[70] = (x[12]);
  assign t[71] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[72] = (x[19]);
  assign t[73] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[74] = (x[25]);
  assign t[75] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[76] = (x[29]);
  assign t[77] = (x[31]);
  assign t[78] = (x[28]);
  assign t[79] = (x[30]);
  assign t[7] = t[11] ? x[15] : t[17];
  assign t[8] = ~(t[16]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[21]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[31]);
  assign t[107] = (x[1]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[40]);
  assign t[111] = (x[0]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[49]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[3]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind141(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[21]);
  assign t[103] = (x[1]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[31]);
  assign t[107] = (x[2]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[40]);
  assign t[111] = (x[3]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[49]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[0]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind146(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[21]);
  assign t[103] = (x[1]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[31]);
  assign t[107] = (x[2]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[40]);
  assign t[111] = (x[3]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[49]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[0]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind151(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [46:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[11]);
  assign t[101] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[102] = (x[33]);
  assign t[103] = (x[6]);
  assign t[104] = (x[12]);
  assign t[105] = (x[40] & ~x[41] & ~x[42] & ~x[43]) | (~x[40] & x[41] & ~x[42] & ~x[43]) | (~x[40] & ~x[41] & x[42] & ~x[43]) | (~x[40] & ~x[41] & ~x[42] & x[43]) | (x[40] & x[41] & x[42] & ~x[43]) | (x[40] & x[41] & ~x[42] & x[43]) | (x[40] & ~x[41] & x[42] & x[43]) | (~x[40] & x[41] & x[42] & x[43]);
  assign t[106] = (x[41]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = t[28] ? t[14] : t[13];
  assign t[12] = ~(t[5] & t[33]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[31] & t[15]);
  assign t[15] = t[8] ? x[29] : t[35];
  assign t[16] = ~(t[17] & t[18]);
  assign t[17] = t[28] ? t[20] : t[19];
  assign t[18] = ~(t[5] & t[32]);
  assign t[19] = ~(t[36]);
  assign t[1] = t[28] ? t[4] : t[3];
  assign t[20] = ~(t[31] & t[21]);
  assign t[21] = t[8] ? x[37] : t[37];
  assign t[22] = ~(t[23] & t[24]);
  assign t[23] = t[28] ? t[26] : t[25];
  assign t[24] = ~(t[5] & t[38]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[31] & t[27]);
  assign t[27] = t[8] ? x[46] : t[40];
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[29]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[30]);
  assign t[40] = (t[53]);
  assign t[41] = t[54] ^ x[2];
  assign t[42] = t[55] ^ x[8];
  assign t[43] = t[56] ^ x[14];
  assign t[44] = t[57] ^ x[17];
  assign t[45] = t[58] ^ x[18];
  assign t[46] = t[59] ^ x[21];
  assign t[47] = t[60] ^ x[22];
  assign t[48] = t[61] ^ x[28];
  assign t[49] = t[62] ^ x[30];
  assign t[4] = ~(t[31] & t[6]);
  assign t[50] = t[63] ^ x[36];
  assign t[51] = t[64] ^ x[38];
  assign t[52] = t[65] ^ x[39];
  assign t[53] = t[66] ^ x[45];
  assign t[54] = (~t[67] & t[68]);
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = (~t[71] & t[72]);
  assign t[57] = (~t[73] & t[74]);
  assign t[58] = (~t[69] & t[75]);
  assign t[59] = (~t[69] & t[76]);
  assign t[5] = ~(t[31] | t[7]);
  assign t[60] = (~t[71] & t[77]);
  assign t[61] = (~t[78] & t[79]);
  assign t[62] = (~t[71] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[69] & t[83]);
  assign t[65] = (~t[71] & t[84]);
  assign t[66] = (~t[85] & t[86]);
  assign t[67] = t[87] ^ x[1];
  assign t[68] = t[88] ^ x[2];
  assign t[69] = t[89] ^ x[7];
  assign t[6] = t[8] ? x[19] : t[32];
  assign t[70] = t[90] ^ x[8];
  assign t[71] = t[91] ^ x[13];
  assign t[72] = t[92] ^ x[14];
  assign t[73] = t[93] ^ x[16];
  assign t[74] = t[94] ^ x[17];
  assign t[75] = t[95] ^ x[18];
  assign t[76] = t[96] ^ x[21];
  assign t[77] = t[97] ^ x[22];
  assign t[78] = t[98] ^ x[27];
  assign t[79] = t[99] ^ x[28];
  assign t[7] = ~(t[28]);
  assign t[80] = t[100] ^ x[30];
  assign t[81] = t[101] ^ x[35];
  assign t[82] = t[102] ^ x[36];
  assign t[83] = t[103] ^ x[38];
  assign t[84] = t[104] ^ x[39];
  assign t[85] = t[105] ^ x[44];
  assign t[86] = t[106] ^ x[45];
  assign t[87] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[0]);
  assign t[89] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[8] = ~(t[9]);
  assign t[90] = (x[3]);
  assign t[91] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[92] = (x[9]);
  assign t[93] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[15]);
  assign t[95] = (x[5]);
  assign t[96] = (x[4]);
  assign t[97] = (x[10]);
  assign t[98] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[99] = (x[25]);
  assign t[9] = ~(x[20]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[22]) | (~t[0] & t[10] & ~t[16] & ~t[22]) | (~t[0] & ~t[10] & t[16] & ~t[22]) | (~t[0] & ~t[10] & ~t[16] & t[22]) | (t[0] & t[10] & t[16] & ~t[22]) | (t[0] & t[10] & ~t[16] & t[22]) | (t[0] & ~t[10] & t[16] & t[22]) | (~t[0] & t[10] & t[16] & t[22]);
endmodule

module R2ind156(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[12]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[5]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[11]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[20]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[4]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[10]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[20]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [20:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[18];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[27] & t[33]);
  assign t[25] = t[34] ^ x[1];
  assign t[26] = t[35] ^ x[2];
  assign t[27] = t[36] ^ x[7];
  assign t[28] = t[37] ^ x[8];
  assign t[29] = t[38] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[39] ^ x[14];
  assign t[31] = t[40] ^ x[16];
  assign t[32] = t[41] ^ x[17];
  assign t[33] = t[42] ^ x[18];
  assign t[34] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[0]);
  assign t[36] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[37] = (x[3]);
  assign t[38] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[5]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[19] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[20]);
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [40:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[9]);
  assign t[10] = ~(x[25]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[37] : t[38];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[40] : t[37];
  assign t[29] = (t[41]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = (t[46]);
  assign t[35] = (t[47]);
  assign t[36] = (t[48]);
  assign t[37] = (t[49]);
  assign t[38] = (t[50]);
  assign t[39] = (t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52]);
  assign t[41] = t[53] ^ x[5];
  assign t[42] = t[54] ^ x[11];
  assign t[43] = t[55] ^ x[14];
  assign t[44] = t[56] ^ x[17];
  assign t[45] = t[57] ^ x[23];
  assign t[46] = t[58] ^ x[26];
  assign t[47] = t[59] ^ x[27];
  assign t[48] = t[60] ^ x[33];
  assign t[49] = t[61] ^ x[35];
  assign t[4] = ~(t[30]);
  assign t[50] = t[62] ^ x[36];
  assign t[51] = t[63] ^ x[38];
  assign t[52] = t[64] ^ x[39];
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[67] & t[68]);
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = (~t[71] & t[72]);
  assign t[57] = (~t[73] & t[74]);
  assign t[58] = (~t[65] & t[75]);
  assign t[59] = (~t[67] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[65] & t[79]);
  assign t[62] = (~t[67] & t[80]);
  assign t[63] = (~t[65] & t[81]);
  assign t[64] = (~t[67] & t[82]);
  assign t[65] = t[83] ^ x[4];
  assign t[66] = t[84] ^ x[5];
  assign t[67] = t[85] ^ x[10];
  assign t[68] = t[86] ^ x[11];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[22];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[32];
  assign t[78] = t[96] ^ x[33];
  assign t[79] = t[97] ^ x[35];
  assign t[7] = ~(t[32]);
  assign t[80] = t[98] ^ x[36];
  assign t[81] = t[99] ^ x[38];
  assign t[82] = t[100] ^ x[39];
  assign t[83] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[84] = (x[0]);
  assign t[85] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[86] = (x[6]);
  assign t[87] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[12]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = (x[15]);
  assign t[91] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[92] = (x[20]);
  assign t[93] = (x[1]);
  assign t[94] = (x[7]);
  assign t[95] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[96] = (x[30]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[3]);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind161(x, y);
 input [20:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[20]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[26] & t[34]);
  assign t[26] = t[35] ^ x[4];
  assign t[27] = t[36] ^ x[5];
  assign t[28] = t[37] ^ x[10];
  assign t[29] = t[38] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[39] ^ x[13];
  assign t[31] = t[40] ^ x[14];
  assign t[32] = t[41] ^ x[16];
  assign t[33] = t[42] ^ x[17];
  assign t[34] = t[43] ^ x[18];
  assign t[35] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[38] = (x[9]);
  assign t[39] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[2]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[19] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [19:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[19]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[5];
  assign t[16] = t[20] ^ x[11];
  assign t[17] = t[21] ^ x[14];
  assign t[18] = t[22] ^ x[17];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[4];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[14];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[17];
  assign t[31] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[32] = (x[2]);
  assign t[33] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[34] = (x[8]);
  assign t[35] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[12]);
  assign t[37] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[15]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[18] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[20]);
  assign t[103] = (x[1]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[30]);
  assign t[107] = (x[2]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[39]);
  assign t[111] = (x[3]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[48]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[0]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind166(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[20]);
  assign t[103] = (x[1]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[30]);
  assign t[107] = (x[2]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[39]);
  assign t[111] = (x[3]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[48]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[0]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind171(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[19]);
  assign t[103] = (x[1]);
  assign t[104] = (x[7]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[29]);
  assign t[107] = (x[2]);
  assign t[108] = (x[8]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(x[25]);
  assign t[110] = (x[38]);
  assign t[111] = (x[3]);
  assign t[112] = (x[9]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[48]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[31] & t[16]);
  assign t[16] = t[9] ? x[34] : t[36];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[37]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[31] & t[22]);
  assign t[22] = t[9] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[31] & t[28]);
  assign t[28] = t[9] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[29]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[30]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[31] & t[8]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[71] & t[81]);
  assign t[63] = (~t[73] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[71] & t[85]);
  assign t[66] = (~t[73] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[71] & t[89]);
  assign t[69] = (~t[73] & t[90]);
  assign t[6] = ~(t[31] | t[7]);
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[4];
  assign t[72] = t[94] ^ x[5];
  assign t[73] = t[95] ^ x[10];
  assign t[74] = t[96] ^ x[11];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[32]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = t[9] ? x[24] : t[33];
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[94] = (x[0]);
  assign t[95] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[96] = (x[6]);
  assign t[97] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[12]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind176(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[20]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[19]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[19]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[0]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[19]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [52:0] x;
 output y;

 wire [115:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[15]);
  assign t[102] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[103] = (x[20]);
  assign t[104] = (x[4]);
  assign t[105] = (x[10]);
  assign t[106] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[107] = (x[29]);
  assign t[108] = (x[5]);
  assign t[109] = (x[11]);
  assign t[10] = ~(t[5] & t[35]);
  assign t[110] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[111] = (x[38]);
  assign t[112] = (x[6]);
  assign t[113] = (x[12]);
  assign t[114] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[115] = (x[47]);
  assign t[11] = ~(t[36]);
  assign t[12] = ~(t[33] & t[13]);
  assign t[13] = t[14] ? x[34] : t[37];
  assign t[14] = ~(t[15]);
  assign t[15] = ~(x[18]);
  assign t[16] = ~(t[17] & t[18]);
  assign t[17] = t[30] ? t[20] : t[19];
  assign t[18] = ~(t[5] & t[38]);
  assign t[19] = ~(t[39]);
  assign t[1] = t[30] ? t[4] : t[3];
  assign t[20] = ~(t[33] & t[21]);
  assign t[21] = t[22] ? x[43] : t[40];
  assign t[22] = ~(t[15]);
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[30] ? t[27] : t[26];
  assign t[25] = ~(t[5] & t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = t[29] ? x[52] : t[43];
  assign t[29] = ~(t[15]);
  assign t[2] = ~(t[5] & t[31]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[32]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = t[58] ^ x[2];
  assign t[45] = t[59] ^ x[8];
  assign t[46] = t[60] ^ x[14];
  assign t[47] = t[61] ^ x[17];
  assign t[48] = t[62] ^ x[24];
  assign t[49] = t[63] ^ x[26];
  assign t[4] = ~(t[33] & t[6]);
  assign t[50] = t[64] ^ x[27];
  assign t[51] = t[65] ^ x[33];
  assign t[52] = t[66] ^ x[35];
  assign t[53] = t[67] ^ x[36];
  assign t[54] = t[68] ^ x[42];
  assign t[55] = t[69] ^ x[44];
  assign t[56] = t[70] ^ x[45];
  assign t[57] = t[71] ^ x[51];
  assign t[58] = (~t[72] & t[73]);
  assign t[59] = (~t[74] & t[75]);
  assign t[5] = ~(t[33] | t[7]);
  assign t[60] = (~t[76] & t[77]);
  assign t[61] = (~t[78] & t[79]);
  assign t[62] = (~t[80] & t[81]);
  assign t[63] = (~t[74] & t[82]);
  assign t[64] = (~t[76] & t[83]);
  assign t[65] = (~t[84] & t[85]);
  assign t[66] = (~t[74] & t[86]);
  assign t[67] = (~t[76] & t[87]);
  assign t[68] = (~t[88] & t[89]);
  assign t[69] = (~t[74] & t[90]);
  assign t[6] = x[18] ? x[25] : t[34];
  assign t[70] = (~t[76] & t[91]);
  assign t[71] = (~t[92] & t[93]);
  assign t[72] = t[94] ^ x[1];
  assign t[73] = t[95] ^ x[2];
  assign t[74] = t[96] ^ x[7];
  assign t[75] = t[97] ^ x[8];
  assign t[76] = t[98] ^ x[13];
  assign t[77] = t[99] ^ x[14];
  assign t[78] = t[100] ^ x[16];
  assign t[79] = t[101] ^ x[17];
  assign t[7] = ~(t[30]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[24];
  assign t[82] = t[104] ^ x[26];
  assign t[83] = t[105] ^ x[27];
  assign t[84] = t[106] ^ x[32];
  assign t[85] = t[107] ^ x[33];
  assign t[86] = t[108] ^ x[35];
  assign t[87] = t[109] ^ x[36];
  assign t[88] = t[110] ^ x[41];
  assign t[89] = t[111] ^ x[42];
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = t[112] ^ x[44];
  assign t[91] = t[113] ^ x[45];
  assign t[92] = t[114] ^ x[50];
  assign t[93] = t[115] ^ x[51];
  assign t[94] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[0]);
  assign t[96] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[97] = (x[3]);
  assign t[98] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[99] = (x[9]);
  assign t[9] = t[30] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[16] & ~t[23]) | (~t[0] & t[8] & ~t[16] & ~t[23]) | (~t[0] & ~t[8] & t[16] & ~t[23]) | (~t[0] & ~t[8] & ~t[16] & t[23]) | (t[0] & t[8] & t[16] & ~t[23]) | (t[0] & t[8] & ~t[16] & t[23]) | (t[0] & ~t[8] & t[16] & t[23]) | (~t[0] & t[8] & t[16] & t[23]);
endmodule

module R2ind181(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[12]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[5]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[11]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[4]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[10]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[10] = ~(t[5] & t[31]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[29] & t[13]);
  assign t[13] = x[18] ? x[29] : t[33];
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = t[26] ? t[18] : t[17];
  assign t[16] = ~(t[5] & t[34]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[29] & t[19]);
  assign t[19] = x[18] ? x[33] : t[36];
  assign t[1] = t[26] ? t[4] : t[3];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[26] ? t[24] : t[23];
  assign t[22] = ~(t[5] & t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] & t[25]);
  assign t[25] = x[18] ? x[36] : t[28];
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = t[52] ^ x[2];
  assign t[3] = ~(t[28]);
  assign t[40] = t[53] ^ x[8];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[24];
  assign t[44] = t[57] ^ x[26];
  assign t[45] = t[58] ^ x[27];
  assign t[46] = t[59] ^ x[28];
  assign t[47] = t[60] ^ x[30];
  assign t[48] = t[61] ^ x[31];
  assign t[49] = t[62] ^ x[32];
  assign t[4] = ~(t[29] & t[6]);
  assign t[50] = t[63] ^ x[34];
  assign t[51] = t[64] ^ x[35];
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = (~t[67] & t[68]);
  assign t[54] = (~t[69] & t[70]);
  assign t[55] = (~t[71] & t[72]);
  assign t[56] = (~t[73] & t[74]);
  assign t[57] = (~t[67] & t[75]);
  assign t[58] = (~t[69] & t[76]);
  assign t[59] = (~t[73] & t[77]);
  assign t[5] = ~(t[29] | t[7]);
  assign t[60] = (~t[67] & t[78]);
  assign t[61] = (~t[69] & t[79]);
  assign t[62] = (~t[73] & t[80]);
  assign t[63] = (~t[67] & t[81]);
  assign t[64] = (~t[69] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[30];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[28];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[31];
  assign t[7] = ~(t[26]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[35];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[21]);
  assign t[96] = (x[5]);
  assign t[97] = (x[11]);
  assign t[98] = (x[22]);
  assign t[99] = (x[6]);
  assign t[9] = t[26] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[14] & ~t[20]) | (~t[0] & t[8] & ~t[14] & ~t[20]) | (~t[0] & ~t[8] & t[14] & ~t[20]) | (~t[0] & ~t[8] & ~t[14] & t[20]) | (t[0] & t[8] & t[14] & ~t[20]) | (t[0] & t[8] & ~t[14] & t[20]) | (t[0] & ~t[8] & t[14] & t[20]) | (~t[0] & t[8] & t[14] & t[20]);
endmodule

module R2ind186(x, y);
 input [20:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[19];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[27] & t[31]);
  assign t[23] = t[32] ^ x[1];
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[39] ^ x[17];
  assign t[31] = t[40] ^ x[19];
  assign t[32] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[0]);
  assign t[34] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[37] = (x[12]);
  assign t[38] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[15]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[20] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[22]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[4]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[10]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[21]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[10] = ~(t[5] & t[31]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[29] & t[13]);
  assign t[13] = x[18] ? x[29] : t[33];
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = t[26] ? t[18] : t[17];
  assign t[16] = ~(t[5] & t[34]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[29] & t[19]);
  assign t[19] = x[18] ? x[33] : t[36];
  assign t[1] = t[26] ? t[4] : t[3];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[26] ? t[24] : t[23];
  assign t[22] = ~(t[5] & t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] & t[25]);
  assign t[25] = x[18] ? x[36] : t[28];
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = t[52] ^ x[2];
  assign t[3] = ~(t[28]);
  assign t[40] = t[53] ^ x[8];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[24];
  assign t[44] = t[57] ^ x[26];
  assign t[45] = t[58] ^ x[27];
  assign t[46] = t[59] ^ x[28];
  assign t[47] = t[60] ^ x[30];
  assign t[48] = t[61] ^ x[31];
  assign t[49] = t[62] ^ x[32];
  assign t[4] = ~(t[29] & t[6]);
  assign t[50] = t[63] ^ x[34];
  assign t[51] = t[64] ^ x[35];
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = (~t[67] & t[68]);
  assign t[54] = (~t[69] & t[70]);
  assign t[55] = (~t[71] & t[72]);
  assign t[56] = (~t[73] & t[74]);
  assign t[57] = (~t[67] & t[75]);
  assign t[58] = (~t[69] & t[76]);
  assign t[59] = (~t[73] & t[77]);
  assign t[5] = ~(t[29] | t[7]);
  assign t[60] = (~t[67] & t[78]);
  assign t[61] = (~t[69] & t[79]);
  assign t[62] = (~t[73] & t[80]);
  assign t[63] = (~t[67] & t[81]);
  assign t[64] = (~t[69] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[30];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[28];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[31];
  assign t[7] = ~(t[26]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[35];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[21]);
  assign t[96] = (x[5]);
  assign t[97] = (x[11]);
  assign t[98] = (x[22]);
  assign t[99] = (x[6]);
  assign t[9] = t[26] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[14] & ~t[20]) | (~t[0] & t[8] & ~t[14] & ~t[20]) | (~t[0] & ~t[8] & t[14] & ~t[20]) | (~t[0] & ~t[8] & ~t[14] & t[20]) | (t[0] & t[8] & t[14] & ~t[20]) | (t[0] & t[8] & ~t[14] & t[20]) | (t[0] & ~t[8] & t[14] & t[20]) | (~t[0] & t[8] & t[14] & t[20]);
endmodule

module R2ind191(x, y);
 input [20:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[19];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[27] & t[31]);
  assign t[23] = t[32] ^ x[1];
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[39] ^ x[17];
  assign t[31] = t[40] ^ x[19];
  assign t[32] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[0]);
  assign t[34] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[37] = (x[12]);
  assign t[38] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[15]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[20] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[22]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[4]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[10]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[21]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind196(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [39:0] x;
 output y;

 wire [109:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[101] = (x[24]);
  assign t[102] = (x[1]);
  assign t[103] = (x[7]);
  assign t[104] = (x[25]);
  assign t[105] = (x[2]);
  assign t[106] = (x[8]);
  assign t[107] = (x[26]);
  assign t[108] = (x[3]);
  assign t[109] = (x[9]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = t[3] ? t[14] : t[13];
  assign t[12] = ~(t[6] & t[34]);
  assign t[13] = ~(t[35]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = x[18] ? x[32] : t[36];
  assign t[16] = ~(t[17] & t[18]);
  assign t[17] = t[3] ? t[20] : t[19];
  assign t[18] = ~(t[6] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[30] & t[21]);
  assign t[21] = x[18] ? x[36] : t[39];
  assign t[22] = ~(t[23] & t[24]);
  assign t[23] = t[3] ? t[26] : t[25];
  assign t[24] = ~(t[6] & t[40]);
  assign t[25] = ~(t[41]);
  assign t[26] = ~(t[30] & t[27]);
  assign t[27] = x[18] ? x[39] : t[29];
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[28]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[11];
  assign t[44] = t[58] ^ x[14];
  assign t[45] = t[59] ^ x[17];
  assign t[46] = t[60] ^ x[22];
  assign t[47] = t[61] ^ x[28];
  assign t[48] = t[62] ^ x[29];
  assign t[49] = t[63] ^ x[30];
  assign t[4] = ~(t[29]);
  assign t[50] = t[64] ^ x[31];
  assign t[51] = t[65] ^ x[33];
  assign t[52] = t[66] ^ x[34];
  assign t[53] = t[67] ^ x[35];
  assign t[54] = t[68] ^ x[37];
  assign t[55] = t[69] ^ x[38];
  assign t[56] = (~t[70] & t[71]);
  assign t[57] = (~t[72] & t[73]);
  assign t[58] = (~t[74] & t[75]);
  assign t[59] = (~t[76] & t[77]);
  assign t[5] = ~(t[30] & t[8]);
  assign t[60] = (~t[78] & t[79]);
  assign t[61] = (~t[80] & t[81]);
  assign t[62] = (~t[70] & t[82]);
  assign t[63] = (~t[72] & t[83]);
  assign t[64] = (~t[80] & t[84]);
  assign t[65] = (~t[70] & t[85]);
  assign t[66] = (~t[72] & t[86]);
  assign t[67] = (~t[80] & t[87]);
  assign t[68] = (~t[70] & t[88]);
  assign t[69] = (~t[72] & t[89]);
  assign t[6] = ~(t[30] | t[7]);
  assign t[70] = t[90] ^ x[4];
  assign t[71] = t[91] ^ x[5];
  assign t[72] = t[92] ^ x[10];
  assign t[73] = t[93] ^ x[11];
  assign t[74] = t[94] ^ x[13];
  assign t[75] = t[95] ^ x[14];
  assign t[76] = t[96] ^ x[16];
  assign t[77] = t[97] ^ x[17];
  assign t[78] = t[98] ^ x[21];
  assign t[79] = t[99] ^ x[22];
  assign t[7] = ~(t[31]);
  assign t[80] = t[100] ^ x[27];
  assign t[81] = t[101] ^ x[28];
  assign t[82] = t[102] ^ x[29];
  assign t[83] = t[103] ^ x[30];
  assign t[84] = t[104] ^ x[31];
  assign t[85] = t[105] ^ x[33];
  assign t[86] = t[106] ^ x[34];
  assign t[87] = t[107] ^ x[35];
  assign t[88] = t[108] ^ x[37];
  assign t[89] = t[109] ^ x[38];
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[90] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[91] = (x[0]);
  assign t[92] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[93] = (x[6]);
  assign t[94] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[12]);
  assign t[96] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[15]);
  assign t[98] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[20]);
  assign t[9] = t[32] ^ t[33];
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[22]) | (~t[0] & t[10] & ~t[16] & ~t[22]) | (~t[0] & ~t[10] & t[16] & ~t[22]) | (~t[0] & ~t[10] & ~t[16] & t[22]) | (t[0] & t[10] & t[16] & ~t[22]) | (t[0] & t[10] & ~t[16] & t[22]) | (t[0] & ~t[10] & t[16] & t[22]) | (~t[0] & t[10] & t[16] & t[22]);
endmodule

module R2ind201(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [28:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[5];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[22];
  assign t[21] = t[27] ^ x[28];
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[38] & t[39]);
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[21];
  assign t[37] = t[49] ^ x[22];
  assign t[38] = t[50] ^ x[27];
  assign t[39] = t[51] ^ x[28];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[6]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[48] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[20]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[51] = (x[24]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [48:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[37];
  assign t[101] = t[127] ^ x[40];
  assign t[102] = t[128] ^ x[41];
  assign t[103] = t[129] ^ x[42];
  assign t[104] = t[130] ^ x[43];
  assign t[105] = t[131] ^ x[44];
  assign t[106] = t[132] ^ x[47];
  assign t[107] = t[133] ^ x[48];
  assign t[108] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[109] = (x[0]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[110] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[111] = (x[6]);
  assign t[112] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[113] = (x[12]);
  assign t[114] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[115] = (x[15]);
  assign t[116] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[20]);
  assign t[118] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[119] = (x[24]);
  assign t[11] = t[3] ? t[14] : t[13];
  assign t[120] = (x[1]);
  assign t[121] = (x[7]);
  assign t[122] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[32]);
  assign t[124] = (x[25]);
  assign t[125] = (x[2]);
  assign t[126] = (x[8]);
  assign t[127] = (x[39] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[39] & 1'b0 & ~1'b0 & ~1'b0) | (~x[39] & ~1'b0 & 1'b0 & ~1'b0) | (~x[39] & ~1'b0 & ~1'b0 & 1'b0) | (x[39] & 1'b0 & 1'b0 & ~1'b0) | (x[39] & 1'b0 & ~1'b0 & 1'b0) | (x[39] & ~1'b0 & 1'b0 & 1'b0) | (~x[39] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[39]);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[6] & t[37]);
  assign t[130] = (x[3]);
  assign t[131] = (x[9]);
  assign t[132] = (x[46] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[46] & 1'b0 & ~1'b0 & ~1'b0) | (~x[46] & ~1'b0 & 1'b0 & ~1'b0) | (~x[46] & ~1'b0 & ~1'b0 & 1'b0) | (x[46] & 1'b0 & 1'b0 & ~1'b0) | (x[46] & 1'b0 & ~1'b0 & 1'b0) | (x[46] & ~1'b0 & 1'b0 & 1'b0) | (~x[46] & 1'b0 & 1'b0 & 1'b0);
  assign t[133] = (x[46]);
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[33] & t[15]);
  assign t[15] = x[18] ? x[31] : t[16];
  assign t[16] = t[39] ^ t[40];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[41]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[42]);
  assign t[21] = ~(t[33] & t[22]);
  assign t[22] = x[18] ? x[38] : t[23];
  assign t[23] = t[43] ^ t[44];
  assign t[24] = ~(t[25] & t[26]);
  assign t[25] = t[3] ? t[28] : t[27];
  assign t[26] = ~(t[6] & t[45]);
  assign t[27] = ~(t[46]);
  assign t[28] = ~(t[33] & t[29]);
  assign t[29] = x[18] ? x[45] : t[30];
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = t[47] ^ t[32];
  assign t[31] = (t[48]);
  assign t[32] = (t[49]);
  assign t[33] = (t[50]);
  assign t[34] = (t[51]);
  assign t[35] = (t[52]);
  assign t[36] = (t[53]);
  assign t[37] = (t[54]);
  assign t[38] = (t[55]);
  assign t[39] = (t[56]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[57]);
  assign t[41] = (t[58]);
  assign t[42] = (t[59]);
  assign t[43] = (t[60]);
  assign t[44] = (t[61]);
  assign t[45] = (t[62]);
  assign t[46] = (t[63]);
  assign t[47] = (t[64]);
  assign t[48] = t[65] ^ x[5];
  assign t[49] = t[66] ^ x[11];
  assign t[4] = ~(t[32]);
  assign t[50] = t[67] ^ x[14];
  assign t[51] = t[68] ^ x[17];
  assign t[52] = t[69] ^ x[22];
  assign t[53] = t[70] ^ x[28];
  assign t[54] = t[71] ^ x[29];
  assign t[55] = t[72] ^ x[30];
  assign t[56] = t[73] ^ x[34];
  assign t[57] = t[74] ^ x[35];
  assign t[58] = t[75] ^ x[36];
  assign t[59] = t[76] ^ x[37];
  assign t[5] = ~(t[33] & t[8]);
  assign t[60] = t[77] ^ x[41];
  assign t[61] = t[78] ^ x[42];
  assign t[62] = t[79] ^ x[43];
  assign t[63] = t[80] ^ x[44];
  assign t[64] = t[81] ^ x[48];
  assign t[65] = (~t[82] & t[83]);
  assign t[66] = (~t[84] & t[85]);
  assign t[67] = (~t[86] & t[87]);
  assign t[68] = (~t[88] & t[89]);
  assign t[69] = (~t[90] & t[91]);
  assign t[6] = ~(t[33] | t[7]);
  assign t[70] = (~t[92] & t[93]);
  assign t[71] = (~t[82] & t[94]);
  assign t[72] = (~t[84] & t[95]);
  assign t[73] = (~t[96] & t[97]);
  assign t[74] = (~t[92] & t[98]);
  assign t[75] = (~t[82] & t[99]);
  assign t[76] = (~t[84] & t[100]);
  assign t[77] = (~t[101] & t[102]);
  assign t[78] = (~t[92] & t[103]);
  assign t[79] = (~t[82] & t[104]);
  assign t[7] = ~(t[34]);
  assign t[80] = (~t[84] & t[105]);
  assign t[81] = (~t[106] & t[107]);
  assign t[82] = t[108] ^ x[4];
  assign t[83] = t[109] ^ x[5];
  assign t[84] = t[110] ^ x[10];
  assign t[85] = t[111] ^ x[11];
  assign t[86] = t[112] ^ x[13];
  assign t[87] = t[113] ^ x[14];
  assign t[88] = t[114] ^ x[16];
  assign t[89] = t[115] ^ x[17];
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[90] = t[116] ^ x[21];
  assign t[91] = t[117] ^ x[22];
  assign t[92] = t[118] ^ x[27];
  assign t[93] = t[119] ^ x[28];
  assign t[94] = t[120] ^ x[29];
  assign t[95] = t[121] ^ x[30];
  assign t[96] = t[122] ^ x[33];
  assign t[97] = t[123] ^ x[34];
  assign t[98] = t[124] ^ x[35];
  assign t[99] = t[125] ^ x[36];
  assign t[9] = t[35] ^ t[36];
  assign y = (t[0] & ~t[10] & ~t[17] & ~t[24]) | (~t[0] & t[10] & ~t[17] & ~t[24]) | (~t[0] & ~t[10] & t[17] & ~t[24]) | (~t[0] & ~t[10] & ~t[17] & t[24]) | (t[0] & t[10] & t[17] & ~t[24]) | (t[0] & t[10] & ~t[17] & t[24]) | (t[0] & ~t[10] & t[17] & t[24]) | (~t[0] & t[10] & t[17] & t[24]);
endmodule

module R2ind206(x, y);
 input [23:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[5];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[22];
  assign t[21] = t[27] ^ x[23];
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[30] & t[38]);
  assign t[28] = t[39] ^ x[4];
  assign t[29] = t[40] ^ x[5];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[41] ^ x[10];
  assign t[31] = t[42] ^ x[11];
  assign t[32] = t[43] ^ x[13];
  assign t[33] = t[44] ^ x[14];
  assign t[34] = t[45] ^ x[16];
  assign t[35] = t[46] ^ x[17];
  assign t[36] = t[47] ^ x[21];
  assign t[37] = t[48] ^ x[22];
  assign t[38] = t[49] ^ x[23];
  assign t[39] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[3]);
  assign t[41] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[44] = (x[12]);
  assign t[45] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[46] = (x[15]);
  assign t[47] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[48] = (x[20]);
  assign t[49] = (x[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [28:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[5];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[22];
  assign t[21] = t[27] ^ x[28];
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[38] & t[39]);
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[21];
  assign t[37] = t[49] ^ x[22];
  assign t[38] = t[50] ^ x[27];
  assign t[39] = t[51] ^ x[28];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[2]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[8]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[48] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[20]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[51] = (x[26]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [28:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[5];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[22];
  assign t[21] = t[27] ^ x[28];
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[38] & t[39]);
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[21];
  assign t[37] = t[49] ^ x[22];
  assign t[38] = t[50] ^ x[27];
  assign t[39] = t[51] ^ x[28];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[48] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[20]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[51] = (x[25]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [28:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[5];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[22];
  assign t[21] = t[27] ^ x[28];
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[38] & t[39]);
  assign t[28] = t[40] ^ x[4];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[21];
  assign t[37] = t[49] ^ x[22];
  assign t[38] = t[50] ^ x[27];
  assign t[39] = t[51] ^ x[28];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[6]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[48] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[20]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[51] = (x[24]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind211(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind216(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind221(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind226(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind231(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [40:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[35]);
  assign t[10] = ~(t[5] & t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[32] & t[13]);
  assign t[13] = t[14] ? x[28] : t[35];
  assign t[14] = ~(t[15]);
  assign t[15] = ~(x[18]);
  assign t[16] = ~(t[17] & t[18]);
  assign t[17] = t[29] ? t[20] : t[19];
  assign t[18] = ~(t[5] & t[36]);
  assign t[19] = ~(t[37]);
  assign t[1] = t[29] ? t[4] : t[3];
  assign t[20] = ~(t[32] & t[21]);
  assign t[21] = t[22] ? x[31] : t[34];
  assign t[22] = ~(t[15]);
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[29] ? t[27] : t[26];
  assign t[25] = ~(t[5] & t[38]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[32] & t[28]);
  assign t[28] = x[18] ? x[40] : t[40];
  assign t[29] = (t[41]);
  assign t[2] = ~(t[5] & t[30]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = (t[46]);
  assign t[35] = (t[47]);
  assign t[36] = (t[48]);
  assign t[37] = (t[49]);
  assign t[38] = (t[50]);
  assign t[39] = (t[51]);
  assign t[3] = ~(t[31]);
  assign t[40] = (t[52]);
  assign t[41] = t[53] ^ x[2];
  assign t[42] = t[54] ^ x[8];
  assign t[43] = t[55] ^ x[14];
  assign t[44] = t[56] ^ x[17];
  assign t[45] = t[57] ^ x[24];
  assign t[46] = t[58] ^ x[26];
  assign t[47] = t[59] ^ x[27];
  assign t[48] = t[60] ^ x[29];
  assign t[49] = t[61] ^ x[30];
  assign t[4] = ~(t[32] & t[6]);
  assign t[50] = t[62] ^ x[32];
  assign t[51] = t[63] ^ x[33];
  assign t[52] = t[64] ^ x[39];
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[67] & t[68]);
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = (~t[71] & t[72]);
  assign t[57] = (~t[73] & t[74]);
  assign t[58] = (~t[67] & t[75]);
  assign t[59] = (~t[69] & t[76]);
  assign t[5] = ~(t[32] | t[7]);
  assign t[60] = (~t[67] & t[77]);
  assign t[61] = (~t[69] & t[78]);
  assign t[62] = (~t[67] & t[79]);
  assign t[63] = (~t[69] & t[80]);
  assign t[64] = (~t[81] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[33];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[29];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[32];
  assign t[7] = ~(t[29]);
  assign t[80] = t[98] ^ x[33];
  assign t[81] = t[99] ^ x[38];
  assign t[82] = t[100] ^ x[39];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[5]);
  assign t[96] = (x[11]);
  assign t[97] = (x[6]);
  assign t[98] = (x[12]);
  assign t[99] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[9] = t[29] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[16] & ~t[23]) | (~t[0] & t[8] & ~t[16] & ~t[23]) | (~t[0] & ~t[8] & t[16] & ~t[23]) | (~t[0] & ~t[8] & ~t[16] & t[23]) | (t[0] & t[8] & t[16] & ~t[23]) | (t[0] & t[8] & ~t[16] & t[23]) | (t[0] & ~t[8] & t[16] & t[23]) | (~t[0] & t[8] & t[16] & t[23]);
endmodule

module R2ind236(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [20:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[18];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[27] & t[33]);
  assign t[25] = t[34] ^ x[1];
  assign t[26] = t[35] ^ x[2];
  assign t[27] = t[36] ^ x[7];
  assign t[28] = t[37] ^ x[8];
  assign t[29] = t[38] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[39] ^ x[14];
  assign t[31] = t[40] ^ x[16];
  assign t[32] = t[41] ^ x[17];
  assign t[33] = t[42] ^ x[18];
  assign t[34] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[0]);
  assign t[36] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[37] = (x[5]);
  assign t[38] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[39] = (x[11]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[4]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[19] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[20]);
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [19:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[2];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[14];
  assign t[17] = t[21] ^ x[17];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = t[30] ^ x[1];
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[7];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[13];
  assign t[27] = t[35] ^ x[14];
  assign t[28] = t[36] ^ x[16];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[0]);
  assign t[32] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[35] = (x[10]);
  assign t[36] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[15]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[18] : t[12];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[19]);
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [52:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[102] = (x[19]);
  assign t[103] = (x[4]);
  assign t[104] = (x[10]);
  assign t[105] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[106] = (x[29]);
  assign t[107] = (x[5]);
  assign t[108] = (x[11]);
  assign t[109] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[110] = (x[38]);
  assign t[111] = (x[6]);
  assign t[112] = (x[12]);
  assign t[113] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[114] = (x[47]);
  assign t[11] = t[29] ? t[14] : t[13];
  assign t[12] = ~(t[5] & t[34]);
  assign t[13] = ~(t[35]);
  assign t[14] = ~(t[32] & t[15]);
  assign t[15] = t[16] ? x[34] : t[36];
  assign t[16] = ~(t[9]);
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[29] ? t[21] : t[20];
  assign t[19] = ~(t[5] & t[37]);
  assign t[1] = t[29] ? t[4] : t[3];
  assign t[20] = ~(t[38]);
  assign t[21] = ~(t[32] & t[22]);
  assign t[22] = x[25] ? x[43] : t[39];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[29] ? t[27] : t[26];
  assign t[25] = ~(t[5] & t[40]);
  assign t[26] = ~(t[41]);
  assign t[27] = ~(t[32] & t[28]);
  assign t[28] = x[25] ? x[52] : t[42];
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[30]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[31]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = t[57] ^ x[2];
  assign t[44] = t[58] ^ x[8];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[23];
  assign t[48] = t[62] ^ x[26];
  assign t[49] = t[63] ^ x[27];
  assign t[4] = ~(t[32] & t[6]);
  assign t[50] = t[64] ^ x[33];
  assign t[51] = t[65] ^ x[35];
  assign t[52] = t[66] ^ x[36];
  assign t[53] = t[67] ^ x[42];
  assign t[54] = t[68] ^ x[44];
  assign t[55] = t[69] ^ x[45];
  assign t[56] = t[70] ^ x[51];
  assign t[57] = (~t[71] & t[72]);
  assign t[58] = (~t[73] & t[74]);
  assign t[59] = (~t[75] & t[76]);
  assign t[5] = ~(t[32] | t[7]);
  assign t[60] = (~t[77] & t[78]);
  assign t[61] = (~t[79] & t[80]);
  assign t[62] = (~t[73] & t[81]);
  assign t[63] = (~t[75] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[73] & t[85]);
  assign t[66] = (~t[75] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[73] & t[89]);
  assign t[69] = (~t[75] & t[90]);
  assign t[6] = t[8] ? x[24] : t[33];
  assign t[70] = (~t[91] & t[92]);
  assign t[71] = t[93] ^ x[1];
  assign t[72] = t[94] ^ x[2];
  assign t[73] = t[95] ^ x[7];
  assign t[74] = t[96] ^ x[8];
  assign t[75] = t[97] ^ x[13];
  assign t[76] = t[98] ^ x[14];
  assign t[77] = t[99] ^ x[16];
  assign t[78] = t[100] ^ x[17];
  assign t[79] = t[101] ^ x[22];
  assign t[7] = ~(t[29]);
  assign t[80] = t[102] ^ x[23];
  assign t[81] = t[103] ^ x[26];
  assign t[82] = t[104] ^ x[27];
  assign t[83] = t[105] ^ x[32];
  assign t[84] = t[106] ^ x[33];
  assign t[85] = t[107] ^ x[35];
  assign t[86] = t[108] ^ x[36];
  assign t[87] = t[109] ^ x[41];
  assign t[88] = t[110] ^ x[42];
  assign t[89] = t[111] ^ x[44];
  assign t[8] = ~(t[9]);
  assign t[90] = t[112] ^ x[45];
  assign t[91] = t[113] ^ x[50];
  assign t[92] = t[114] ^ x[51];
  assign t[93] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[0]);
  assign t[95] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[96] = (x[3]);
  assign t[97] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[98] = (x[9]);
  assign t[99] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(x[25]);
  assign y = (t[0] & ~t[10] & ~t[17] & ~t[23]) | (~t[0] & t[10] & ~t[17] & ~t[23]) | (~t[0] & ~t[10] & t[17] & ~t[23]) | (~t[0] & ~t[10] & ~t[17] & t[23]) | (t[0] & t[10] & t[17] & ~t[23]) | (t[0] & t[10] & ~t[17] & t[23]) | (t[0] & ~t[10] & t[17] & t[23]) | (~t[0] & t[10] & t[17] & t[23]);
endmodule

module R2ind241(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[4]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[10]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [25:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[17];
  assign t[19] = t[24] ^ x[23];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[0]);
  assign t[37] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[38] = (x[3]);
  assign t[39] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[9]);
  assign t[41] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[42] = (x[15]);
  assign t[43] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[44] = (x[19]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[24] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[25]);
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [52:0] x;
 output y;

 wire [116:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[101] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[15]);
  assign t[103] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[104] = (x[19]);
  assign t[105] = (x[1]);
  assign t[106] = (x[7]);
  assign t[107] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[108] = (x[28]);
  assign t[109] = (x[2]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[110] = (x[8]);
  assign t[111] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[112] = (x[37]);
  assign t[113] = (x[3]);
  assign t[114] = (x[9]);
  assign t[115] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[116] = (x[49]);
  assign t[11] = ~(t[6] & t[36]);
  assign t[12] = ~(t[37]);
  assign t[13] = ~(t[33] & t[14]);
  assign t[14] = t[15] ? x[34] : t[38];
  assign t[15] = ~(t[16]);
  assign t[16] = ~(x[18]);
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[39]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[40]);
  assign t[21] = ~(t[33] & t[22]);
  assign t[22] = t[23] ? x[43] : t[41];
  assign t[23] = ~(t[16]);
  assign t[24] = ~(t[25] & t[26]);
  assign t[25] = t[3] ? t[28] : t[27];
  assign t[26] = ~(t[6] & t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[33] & t[29]);
  assign t[29] = t[30] ? x[52] : t[44];
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[16]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = t[59] ^ x[5];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[14];
  assign t[48] = t[62] ^ x[17];
  assign t[49] = t[63] ^ x[24];
  assign t[4] = ~(t[32]);
  assign t[50] = t[64] ^ x[26];
  assign t[51] = t[65] ^ x[27];
  assign t[52] = t[66] ^ x[33];
  assign t[53] = t[67] ^ x[35];
  assign t[54] = t[68] ^ x[36];
  assign t[55] = t[69] ^ x[42];
  assign t[56] = t[70] ^ x[44];
  assign t[57] = t[71] ^ x[45];
  assign t[58] = t[72] ^ x[51];
  assign t[59] = (~t[73] & t[74]);
  assign t[5] = ~(t[33] & t[8]);
  assign t[60] = (~t[75] & t[76]);
  assign t[61] = (~t[77] & t[78]);
  assign t[62] = (~t[79] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[73] & t[83]);
  assign t[65] = (~t[75] & t[84]);
  assign t[66] = (~t[85] & t[86]);
  assign t[67] = (~t[73] & t[87]);
  assign t[68] = (~t[75] & t[88]);
  assign t[69] = (~t[89] & t[90]);
  assign t[6] = ~(t[33] | t[7]);
  assign t[70] = (~t[73] & t[91]);
  assign t[71] = (~t[75] & t[92]);
  assign t[72] = (~t[93] & t[94]);
  assign t[73] = t[95] ^ x[4];
  assign t[74] = t[96] ^ x[5];
  assign t[75] = t[97] ^ x[10];
  assign t[76] = t[98] ^ x[11];
  assign t[77] = t[99] ^ x[13];
  assign t[78] = t[100] ^ x[14];
  assign t[79] = t[101] ^ x[16];
  assign t[7] = ~(t[34]);
  assign t[80] = t[102] ^ x[17];
  assign t[81] = t[103] ^ x[23];
  assign t[82] = t[104] ^ x[24];
  assign t[83] = t[105] ^ x[26];
  assign t[84] = t[106] ^ x[27];
  assign t[85] = t[107] ^ x[32];
  assign t[86] = t[108] ^ x[33];
  assign t[87] = t[109] ^ x[35];
  assign t[88] = t[110] ^ x[36];
  assign t[89] = t[111] ^ x[41];
  assign t[8] = x[18] ? x[25] : t[35];
  assign t[90] = t[112] ^ x[42];
  assign t[91] = t[113] ^ x[44];
  assign t[92] = t[114] ^ x[45];
  assign t[93] = t[115] ^ x[50];
  assign t[94] = t[116] ^ x[51];
  assign t[95] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[96] = (x[0]);
  assign t[97] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[98] = (x[6]);
  assign t[99] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[17] & ~t[24]) | (~t[0] & t[9] & ~t[17] & ~t[24]) | (~t[0] & ~t[9] & t[17] & ~t[24]) | (~t[0] & ~t[9] & ~t[17] & t[24]) | (t[0] & t[9] & t[17] & ~t[24]) | (t[0] & t[9] & ~t[17] & t[24]) | (t[0] & ~t[9] & t[17] & t[24]) | (~t[0] & t[9] & t[17] & t[24]);
endmodule

module R2ind246(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[21]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[18]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[7]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[18]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [52:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[1]);
  assign t[102] = (x[7]);
  assign t[103] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[104] = (x[28]);
  assign t[105] = (x[2]);
  assign t[106] = (x[8]);
  assign t[107] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[108] = (x[37]);
  assign t[109] = (x[3]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[110] = (x[9]);
  assign t[111] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[112] = (x[46]);
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[34] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[43] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[52] : t[40];
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = t[55] ^ x[5];
  assign t[42] = t[56] ^ x[11];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[24];
  assign t[46] = t[60] ^ x[26];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[33];
  assign t[49] = t[63] ^ x[35];
  assign t[4] = ~(t[28]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[42];
  assign t[52] = t[66] ^ x[44];
  assign t[53] = t[67] ^ x[45];
  assign t[54] = t[68] ^ x[51];
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = (~t[71] & t[72]);
  assign t[57] = (~t[73] & t[74]);
  assign t[58] = (~t[75] & t[76]);
  assign t[59] = (~t[77] & t[78]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[69] & t[79]);
  assign t[61] = (~t[71] & t[80]);
  assign t[62] = (~t[81] & t[82]);
  assign t[63] = (~t[69] & t[83]);
  assign t[64] = (~t[71] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[69] & t[87]);
  assign t[67] = (~t[71] & t[88]);
  assign t[68] = (~t[89] & t[90]);
  assign t[69] = t[91] ^ x[4];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[92] ^ x[5];
  assign t[71] = t[93] ^ x[10];
  assign t[72] = t[94] ^ x[11];
  assign t[73] = t[95] ^ x[13];
  assign t[74] = t[96] ^ x[14];
  assign t[75] = t[97] ^ x[16];
  assign t[76] = t[98] ^ x[17];
  assign t[77] = t[99] ^ x[23];
  assign t[78] = t[100] ^ x[24];
  assign t[79] = t[101] ^ x[26];
  assign t[7] = ~(t[30]);
  assign t[80] = t[102] ^ x[27];
  assign t[81] = t[103] ^ x[32];
  assign t[82] = t[104] ^ x[33];
  assign t[83] = t[105] ^ x[35];
  assign t[84] = t[106] ^ x[36];
  assign t[85] = t[107] ^ x[41];
  assign t[86] = t[108] ^ x[42];
  assign t[87] = t[109] ^ x[44];
  assign t[88] = t[110] ^ x[45];
  assign t[89] = t[111] ^ x[50];
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = t[112] ^ x[51];
  assign t[91] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[92] = (x[0]);
  assign t[93] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[94] = (x[6]);
  assign t[95] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[12]);
  assign t[97] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[15]);
  assign t[99] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind251(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[9]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [52:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[1]);
  assign t[102] = (x[7]);
  assign t[103] = (x[28] & ~x[29] & ~x[30] & ~x[31]) | (~x[28] & x[29] & ~x[30] & ~x[31]) | (~x[28] & ~x[29] & x[30] & ~x[31]) | (~x[28] & ~x[29] & ~x[30] & x[31]) | (x[28] & x[29] & x[30] & ~x[31]) | (x[28] & x[29] & ~x[30] & x[31]) | (x[28] & ~x[29] & x[30] & x[31]) | (~x[28] & x[29] & x[30] & x[31]);
  assign t[104] = (x[28]);
  assign t[105] = (x[2]);
  assign t[106] = (x[8]);
  assign t[107] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[108] = (x[37]);
  assign t[109] = (x[3]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[110] = (x[9]);
  assign t[111] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[112] = (x[46]);
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[34] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[43] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[52] : t[40];
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[54]);
  assign t[41] = t[55] ^ x[5];
  assign t[42] = t[56] ^ x[11];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[24];
  assign t[46] = t[60] ^ x[26];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[33];
  assign t[49] = t[63] ^ x[35];
  assign t[4] = ~(t[28]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[42];
  assign t[52] = t[66] ^ x[44];
  assign t[53] = t[67] ^ x[45];
  assign t[54] = t[68] ^ x[51];
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = (~t[71] & t[72]);
  assign t[57] = (~t[73] & t[74]);
  assign t[58] = (~t[75] & t[76]);
  assign t[59] = (~t[77] & t[78]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[69] & t[79]);
  assign t[61] = (~t[71] & t[80]);
  assign t[62] = (~t[81] & t[82]);
  assign t[63] = (~t[69] & t[83]);
  assign t[64] = (~t[71] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[69] & t[87]);
  assign t[67] = (~t[71] & t[88]);
  assign t[68] = (~t[89] & t[90]);
  assign t[69] = t[91] ^ x[4];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[92] ^ x[5];
  assign t[71] = t[93] ^ x[10];
  assign t[72] = t[94] ^ x[11];
  assign t[73] = t[95] ^ x[13];
  assign t[74] = t[96] ^ x[14];
  assign t[75] = t[97] ^ x[16];
  assign t[76] = t[98] ^ x[17];
  assign t[77] = t[99] ^ x[23];
  assign t[78] = t[100] ^ x[24];
  assign t[79] = t[101] ^ x[26];
  assign t[7] = ~(t[30]);
  assign t[80] = t[102] ^ x[27];
  assign t[81] = t[103] ^ x[32];
  assign t[82] = t[104] ^ x[33];
  assign t[83] = t[105] ^ x[35];
  assign t[84] = t[106] ^ x[36];
  assign t[85] = t[107] ^ x[41];
  assign t[86] = t[108] ^ x[42];
  assign t[87] = t[109] ^ x[44];
  assign t[88] = t[110] ^ x[45];
  assign t[89] = t[111] ^ x[50];
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = t[112] ^ x[51];
  assign t[91] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[92] = (x[0]);
  assign t[93] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[94] = (x[6]);
  assign t[95] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[12]);
  assign t[97] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[15]);
  assign t[99] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind256(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[9]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[19]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [40:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[101] = (x[34]);
  assign t[10] = ~(x[19]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = t[3] ? t[15] : t[14];
  assign t[13] = ~(t[6] & t[34]);
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[32] & t[16]);
  assign t[16] = x[19] ? x[22] : t[30];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = t[3] ? t[21] : t[20];
  assign t[19] = ~(t[6] & t[36]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[37]);
  assign t[21] = ~(t[32] & t[22]);
  assign t[22] = t[9] ? x[31] : t[38];
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = t[3] ? t[27] : t[26];
  assign t[25] = ~(t[6] & t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[32] & t[28]);
  assign t[28] = t[29] ? x[40] : t[41];
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = (t[46]);
  assign t[35] = (t[47]);
  assign t[36] = (t[48]);
  assign t[37] = (t[49]);
  assign t[38] = (t[50]);
  assign t[39] = (t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52]);
  assign t[41] = (t[53]);
  assign t[42] = t[54] ^ x[5];
  assign t[43] = t[55] ^ x[11];
  assign t[44] = t[56] ^ x[14];
  assign t[45] = t[57] ^ x[17];
  assign t[46] = t[58] ^ x[20];
  assign t[47] = t[59] ^ x[21];
  assign t[48] = t[60] ^ x[23];
  assign t[49] = t[61] ^ x[24];
  assign t[4] = ~(t[31]);
  assign t[50] = t[62] ^ x[30];
  assign t[51] = t[63] ^ x[32];
  assign t[52] = t[64] ^ x[33];
  assign t[53] = t[65] ^ x[39];
  assign t[54] = (~t[66] & t[67]);
  assign t[55] = (~t[68] & t[69]);
  assign t[56] = (~t[70] & t[71]);
  assign t[57] = (~t[72] & t[73]);
  assign t[58] = (~t[66] & t[74]);
  assign t[59] = (~t[68] & t[75]);
  assign t[5] = ~(t[32] & t[8]);
  assign t[60] = (~t[66] & t[76]);
  assign t[61] = (~t[68] & t[77]);
  assign t[62] = (~t[78] & t[79]);
  assign t[63] = (~t[66] & t[80]);
  assign t[64] = (~t[68] & t[81]);
  assign t[65] = (~t[82] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[32] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[20];
  assign t[75] = t[93] ^ x[21];
  assign t[76] = t[94] ^ x[23];
  assign t[77] = t[95] ^ x[24];
  assign t[78] = t[96] ^ x[29];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[33]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[33];
  assign t[82] = t[100] ^ x[38];
  assign t[83] = t[101] ^ x[39];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = t[9] ? x[18] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[1]);
  assign t[93] = (x[7]);
  assign t[94] = (x[2]);
  assign t[95] = (x[8]);
  assign t[96] = (x[25] & ~x[26] & ~x[27] & ~x[28]) | (~x[25] & x[26] & ~x[27] & ~x[28]) | (~x[25] & ~x[26] & x[27] & ~x[28]) | (~x[25] & ~x[26] & ~x[27] & x[28]) | (x[25] & x[26] & x[27] & ~x[28]) | (x[25] & x[26] & ~x[27] & x[28]) | (x[25] & ~x[26] & x[27] & x[28]) | (~x[25] & x[26] & x[27] & x[28]);
  assign t[97] = (x[25]);
  assign t[98] = (x[3]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[11] & ~t[17] & ~t[23]) | (~t[0] & t[11] & ~t[17] & ~t[23]) | (~t[0] & ~t[11] & t[17] & ~t[23]) | (~t[0] & ~t[11] & ~t[17] & t[23]) | (t[0] & t[11] & t[17] & ~t[23]) | (t[0] & t[11] & ~t[17] & t[23]) | (t[0] & ~t[11] & t[17] & t[23]) | (~t[0] & t[11] & t[17] & t[23]);
endmodule

module R2ind261(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[18]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[25]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[14];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[23];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[13];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[17];
  assign t[34] = t[44] ^ x[22];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[2]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[8]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[12]);
  assign t[42] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[15]);
  assign t[44] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[45] = (x[18]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[24] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[24] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[7]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[0]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [19:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[19]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[5];
  assign t[16] = t[20] ^ x[11];
  assign t[17] = t[21] ^ x[14];
  assign t[18] = t[22] ^ x[17];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[4];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[13];
  assign t[28] = t[36] ^ x[14];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[17];
  assign t[31] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[32] = (x[0]);
  assign t[33] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[34] = (x[6]);
  assign t[35] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[12]);
  assign t[37] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[15]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[18] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind266(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind271(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[10] = ~(t[5] & t[31]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[29] & t[13]);
  assign t[13] = x[18] ? x[29] : t[33];
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = t[26] ? t[18] : t[17];
  assign t[16] = ~(t[5] & t[34]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[29] & t[19]);
  assign t[19] = x[18] ? x[33] : t[36];
  assign t[1] = t[26] ? t[4] : t[3];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[26] ? t[24] : t[23];
  assign t[22] = ~(t[5] & t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] & t[25]);
  assign t[25] = x[18] ? x[36] : t[28];
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = t[52] ^ x[2];
  assign t[3] = ~(t[28]);
  assign t[40] = t[53] ^ x[8];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[24];
  assign t[44] = t[57] ^ x[26];
  assign t[45] = t[58] ^ x[27];
  assign t[46] = t[59] ^ x[28];
  assign t[47] = t[60] ^ x[30];
  assign t[48] = t[61] ^ x[31];
  assign t[49] = t[62] ^ x[32];
  assign t[4] = ~(t[29] & t[6]);
  assign t[50] = t[63] ^ x[34];
  assign t[51] = t[64] ^ x[35];
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = (~t[67] & t[68]);
  assign t[54] = (~t[69] & t[70]);
  assign t[55] = (~t[71] & t[72]);
  assign t[56] = (~t[73] & t[74]);
  assign t[57] = (~t[67] & t[75]);
  assign t[58] = (~t[69] & t[76]);
  assign t[59] = (~t[73] & t[77]);
  assign t[5] = ~(t[29] | t[7]);
  assign t[60] = (~t[67] & t[78]);
  assign t[61] = (~t[69] & t[79]);
  assign t[62] = (~t[73] & t[80]);
  assign t[63] = (~t[67] & t[81]);
  assign t[64] = (~t[69] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[30];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[28];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[31];
  assign t[7] = ~(t[26]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[35];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[21]);
  assign t[96] = (x[5]);
  assign t[97] = (x[11]);
  assign t[98] = (x[22]);
  assign t[99] = (x[6]);
  assign t[9] = t[26] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[14] & ~t[20]) | (~t[0] & t[8] & ~t[14] & ~t[20]) | (~t[0] & ~t[8] & t[14] & ~t[20]) | (~t[0] & ~t[8] & ~t[14] & t[20]) | (t[0] & t[8] & t[14] & ~t[20]) | (t[0] & t[8] & ~t[14] & t[20]) | (t[0] & ~t[8] & t[14] & t[20]) | (~t[0] & t[8] & t[14] & t[20]);
endmodule

module R2ind276(x, y);
 input [20:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[19];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[27] & t[31]);
  assign t[23] = t[32] ^ x[1];
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[39] ^ x[17];
  assign t[31] = t[40] ^ x[19];
  assign t[32] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[0]);
  assign t[34] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[37] = (x[12]);
  assign t[38] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[15]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[20] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[22]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[4]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[10]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[21]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[10] = ~(t[5] & t[31]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[29] & t[13]);
  assign t[13] = x[18] ? x[29] : t[33];
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = t[26] ? t[18] : t[17];
  assign t[16] = ~(t[5] & t[34]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[29] & t[19]);
  assign t[19] = x[18] ? x[33] : t[36];
  assign t[1] = t[26] ? t[4] : t[3];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[26] ? t[24] : t[23];
  assign t[22] = ~(t[5] & t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] & t[25]);
  assign t[25] = x[18] ? x[36] : t[28];
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = t[52] ^ x[2];
  assign t[3] = ~(t[28]);
  assign t[40] = t[53] ^ x[8];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[24];
  assign t[44] = t[57] ^ x[26];
  assign t[45] = t[58] ^ x[27];
  assign t[46] = t[59] ^ x[28];
  assign t[47] = t[60] ^ x[30];
  assign t[48] = t[61] ^ x[31];
  assign t[49] = t[62] ^ x[32];
  assign t[4] = ~(t[29] & t[6]);
  assign t[50] = t[63] ^ x[34];
  assign t[51] = t[64] ^ x[35];
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = (~t[67] & t[68]);
  assign t[54] = (~t[69] & t[70]);
  assign t[55] = (~t[71] & t[72]);
  assign t[56] = (~t[73] & t[74]);
  assign t[57] = (~t[67] & t[75]);
  assign t[58] = (~t[69] & t[76]);
  assign t[59] = (~t[73] & t[77]);
  assign t[5] = ~(t[29] | t[7]);
  assign t[60] = (~t[67] & t[78]);
  assign t[61] = (~t[69] & t[79]);
  assign t[62] = (~t[73] & t[80]);
  assign t[63] = (~t[67] & t[81]);
  assign t[64] = (~t[69] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[30];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[28];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[31];
  assign t[7] = ~(t[26]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[35];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[21]);
  assign t[96] = (x[5]);
  assign t[97] = (x[11]);
  assign t[98] = (x[22]);
  assign t[99] = (x[6]);
  assign t[9] = t[26] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[14] & ~t[20]) | (~t[0] & t[8] & ~t[14] & ~t[20]) | (~t[0] & ~t[8] & t[14] & ~t[20]) | (~t[0] & ~t[8] & ~t[14] & t[20]) | (t[0] & t[8] & t[14] & ~t[20]) | (t[0] & t[8] & ~t[14] & t[20]) | (t[0] & ~t[8] & t[14] & t[20]) | (~t[0] & t[8] & t[14] & t[20]);
endmodule

module R2ind281(x, y);
 input [20:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[19];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[27] & t[31]);
  assign t[23] = t[32] ^ x[1];
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[39] ^ x[17];
  assign t[31] = t[40] ^ x[19];
  assign t[32] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[0]);
  assign t[34] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[37] = (x[12]);
  assign t[38] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[15]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[20] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[22]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[4]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[10]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[21]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[12]);
  assign t[10] = ~(t[5] & t[31]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[29] & t[13]);
  assign t[13] = x[18] ? x[29] : t[33];
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = t[26] ? t[18] : t[17];
  assign t[16] = ~(t[5] & t[34]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[29] & t[19]);
  assign t[19] = x[18] ? x[33] : t[36];
  assign t[1] = t[26] ? t[4] : t[3];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[26] ? t[24] : t[23];
  assign t[22] = ~(t[5] & t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] & t[25]);
  assign t[25] = x[18] ? x[36] : t[28];
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[5] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = t[52] ^ x[2];
  assign t[3] = ~(t[28]);
  assign t[40] = t[53] ^ x[8];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[24];
  assign t[44] = t[57] ^ x[26];
  assign t[45] = t[58] ^ x[27];
  assign t[46] = t[59] ^ x[28];
  assign t[47] = t[60] ^ x[30];
  assign t[48] = t[61] ^ x[31];
  assign t[49] = t[62] ^ x[32];
  assign t[4] = ~(t[29] & t[6]);
  assign t[50] = t[63] ^ x[34];
  assign t[51] = t[64] ^ x[35];
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = (~t[67] & t[68]);
  assign t[54] = (~t[69] & t[70]);
  assign t[55] = (~t[71] & t[72]);
  assign t[56] = (~t[73] & t[74]);
  assign t[57] = (~t[67] & t[75]);
  assign t[58] = (~t[69] & t[76]);
  assign t[59] = (~t[73] & t[77]);
  assign t[5] = ~(t[29] | t[7]);
  assign t[60] = (~t[67] & t[78]);
  assign t[61] = (~t[69] & t[79]);
  assign t[62] = (~t[73] & t[80]);
  assign t[63] = (~t[67] & t[81]);
  assign t[64] = (~t[69] & t[82]);
  assign t[65] = t[83] ^ x[1];
  assign t[66] = t[84] ^ x[2];
  assign t[67] = t[85] ^ x[7];
  assign t[68] = t[86] ^ x[8];
  assign t[69] = t[87] ^ x[13];
  assign t[6] = x[18] ? x[25] : t[30];
  assign t[70] = t[88] ^ x[14];
  assign t[71] = t[89] ^ x[16];
  assign t[72] = t[90] ^ x[17];
  assign t[73] = t[91] ^ x[23];
  assign t[74] = t[92] ^ x[24];
  assign t[75] = t[93] ^ x[26];
  assign t[76] = t[94] ^ x[27];
  assign t[77] = t[95] ^ x[28];
  assign t[78] = t[96] ^ x[30];
  assign t[79] = t[97] ^ x[31];
  assign t[7] = ~(t[26]);
  assign t[80] = t[98] ^ x[32];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[35];
  assign t[83] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[0]);
  assign t[85] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[86] = (x[3]);
  assign t[87] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[88] = (x[9]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] & t[10]);
  assign t[90] = (x[15]);
  assign t[91] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[92] = (x[20]);
  assign t[93] = (x[4]);
  assign t[94] = (x[10]);
  assign t[95] = (x[21]);
  assign t[96] = (x[5]);
  assign t[97] = (x[11]);
  assign t[98] = (x[22]);
  assign t[99] = (x[6]);
  assign t[9] = t[26] ? t[12] : t[11];
  assign y = (t[0] & ~t[8] & ~t[14] & ~t[20]) | (~t[0] & t[8] & ~t[14] & ~t[20]) | (~t[0] & ~t[8] & t[14] & ~t[20]) | (~t[0] & ~t[8] & ~t[14] & t[20]) | (t[0] & t[8] & t[14] & ~t[20]) | (t[0] & t[8] & ~t[14] & t[20]) | (t[0] & ~t[8] & t[14] & t[20]) | (~t[0] & t[8] & t[14] & t[20]);
endmodule

module R2ind286(x, y);
 input [20:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[19];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[27] & t[31]);
  assign t[23] = t[32] ^ x[1];
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[39] ^ x[17];
  assign t[31] = t[40] ^ x[19];
  assign t[32] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[0]);
  assign t[34] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[37] = (x[12]);
  assign t[38] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[15]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[20] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[5]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[22]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[4]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[10]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[21]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[8];
  assign t[15] = t[20] ^ x[14];
  assign t[16] = t[21] ^ x[17];
  assign t[17] = t[22] ^ x[24];
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[25] & t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (~t[27] & t[28]);
  assign t[21] = (~t[29] & t[30]);
  assign t[22] = (~t[31] & t[32]);
  assign t[23] = t[33] ^ x[1];
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[7];
  assign t[26] = t[36] ^ x[8];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[14];
  assign t[29] = t[39] ^ x[16];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[23];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[0]);
  assign t[35] = (x[3] & ~x[4] & ~x[5] & ~x[6]) | (~x[3] & x[4] & ~x[5] & ~x[6]) | (~x[3] & ~x[4] & x[5] & ~x[6]) | (~x[3] & ~x[4] & ~x[5] & x[6]) | (x[3] & x[4] & x[5] & ~x[6]) | (x[3] & x[4] & ~x[5] & x[6]) | (x[3] & ~x[4] & x[5] & x[6]) | (~x[3] & x[4] & x[5] & x[6]);
  assign t[36] = (x[3]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[9]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[15]);
  assign t[41] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[42] = (x[20]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[18] ? x[25] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind291(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind296(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind301(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [36:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[10] = t[3] ? t[13] : t[12];
  assign t[11] = ~(t[6] & t[32]);
  assign t[12] = ~(t[33]);
  assign t[13] = ~(t[29] & t[14]);
  assign t[14] = x[18] ? x[29] : t[34];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = t[3] ? t[19] : t[18];
  assign t[17] = ~(t[6] & t[35]);
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[29] & t[20]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = x[18] ? x[33] : t[37];
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = t[3] ? t[25] : t[24];
  assign t[23] = ~(t[6] & t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[29] & t[26]);
  assign t[26] = x[18] ? x[36] : t[28];
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[6] & t[27]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[5];
  assign t[41] = t[54] ^ x[11];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[17];
  assign t[44] = t[57] ^ x[24];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[27];
  assign t[47] = t[60] ^ x[28];
  assign t[48] = t[61] ^ x[30];
  assign t[49] = t[62] ^ x[31];
  assign t[4] = ~(t[28]);
  assign t[50] = t[63] ^ x[32];
  assign t[51] = t[64] ^ x[34];
  assign t[52] = t[65] ^ x[35];
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[72] & t[73]);
  assign t[57] = (~t[74] & t[75]);
  assign t[58] = (~t[66] & t[76]);
  assign t[59] = (~t[68] & t[77]);
  assign t[5] = ~(t[29] & t[8]);
  assign t[60] = (~t[74] & t[78]);
  assign t[61] = (~t[66] & t[79]);
  assign t[62] = (~t[68] & t[80]);
  assign t[63] = (~t[74] & t[81]);
  assign t[64] = (~t[66] & t[82]);
  assign t[65] = (~t[68] & t[83]);
  assign t[66] = t[84] ^ x[4];
  assign t[67] = t[85] ^ x[5];
  assign t[68] = t[86] ^ x[10];
  assign t[69] = t[87] ^ x[11];
  assign t[6] = ~(t[29] | t[7]);
  assign t[70] = t[88] ^ x[13];
  assign t[71] = t[89] ^ x[14];
  assign t[72] = t[90] ^ x[16];
  assign t[73] = t[91] ^ x[17];
  assign t[74] = t[92] ^ x[23];
  assign t[75] = t[93] ^ x[24];
  assign t[76] = t[94] ^ x[26];
  assign t[77] = t[95] ^ x[27];
  assign t[78] = t[96] ^ x[28];
  assign t[79] = t[97] ^ x[30];
  assign t[7] = ~(t[30]);
  assign t[80] = t[98] ^ x[31];
  assign t[81] = t[99] ^ x[32];
  assign t[82] = t[100] ^ x[34];
  assign t[83] = t[101] ^ x[35];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[87] = (x[6]);
  assign t[88] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[12]);
  assign t[8] = x[18] ? x[25] : t[31];
  assign t[90] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[15]);
  assign t[92] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[93] = (x[20]);
  assign t[94] = (x[1]);
  assign t[95] = (x[7]);
  assign t[96] = (x[21]);
  assign t[97] = (x[2]);
  assign t[98] = (x[8]);
  assign t[99] = (x[22]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[9] & ~t[15] & ~t[21]) | (~t[0] & t[9] & ~t[15] & ~t[21]) | (~t[0] & ~t[9] & t[15] & ~t[21]) | (~t[0] & ~t[9] & ~t[15] & t[21]) | (t[0] & t[9] & t[15] & ~t[21]) | (t[0] & t[9] & ~t[15] & t[21]) | (t[0] & ~t[9] & t[15] & t[21]) | (~t[0] & t[9] & t[15] & t[21]);
endmodule

module R2ind306(x, y);
 input [20:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[19];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[26] & t[32]);
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[39] ^ x[16];
  assign t[31] = t[40] ^ x[17];
  assign t[32] = t[41] ^ x[19];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[36] = (x[9]);
  assign t[37] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[12]);
  assign t[39] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15]);
  assign t[41] = (x[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[20] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[2]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[8]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[22]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[7]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[21]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [25:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[14];
  assign t[17] = t[22] ^ x[17];
  assign t[18] = t[23] ^ x[24];
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = (~t[30] & t[31]);
  assign t[23] = (~t[32] & t[33]);
  assign t[24] = t[34] ^ x[4];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[13];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[17];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[0]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[12]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[15]);
  assign t[42] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[43] = (x[20]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[18] ? x[25] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [37:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[119] ^ x[16];
  assign t[101] = t[120] ^ x[17];
  assign t[102] = t[121] ^ x[24];
  assign t[103] = t[122] ^ x[25];
  assign t[104] = t[123] ^ x[26];
  assign t[105] = t[124] ^ x[27];
  assign t[106] = t[125] ^ x[28];
  assign t[107] = t[126] ^ x[29];
  assign t[108] = t[127] ^ x[30];
  assign t[109] = t[128] ^ x[32];
  assign t[10] = t[56] ? t[13] : t[12];
  assign t[110] = t[129] ^ x[33];
  assign t[111] = t[130] ^ x[35];
  assign t[112] = t[131] ^ x[36];
  assign t[113] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[114] = (x[0]);
  assign t[115] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[116] = (x[6]);
  assign t[117] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[12]);
  assign t[119] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[14] & t[15]);
  assign t[120] = (x[15]);
  assign t[121] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[122] = (x[23]);
  assign t[123] = (x[21]);
  assign t[124] = (x[20]);
  assign t[125] = (x[22]);
  assign t[126] = (x[1]);
  assign t[127] = (x[7]);
  assign t[128] = (x[2]);
  assign t[129] = (x[8]);
  assign t[12] = ~(t[57] & t[16]);
  assign t[130] = (x[3]);
  assign t[131] = (x[9]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[56] | t[58]);
  assign t[15] = ~(t[57]);
  assign t[16] = ~(t[19] & t[17]);
  assign t[17] = ~(t[59]);
  assign t[18] = ~(t[19] & t[15]);
  assign t[19] = ~(t[58]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = t[3] ? t[24] : t[23];
  assign t[22] = ~(t[6] & t[60]);
  assign t[23] = ~(t[61]);
  assign t[24] = ~(t[54] & t[25]);
  assign t[25] = x[18] ? x[31] : t[26];
  assign t[26] = ~(t[27] & t[28]);
  assign t[27] = ~(t[29] & t[12]);
  assign t[28] = ~(t[30] & t[31]);
  assign t[29] = ~(t[59] | t[32]);
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[14] | t[17]);
  assign t[31] = t[56] ? t[12] : t[57];
  assign t[32] = ~(t[33] | t[18]);
  assign t[33] = ~(t[56]);
  assign t[34] = ~(t[35] & t[36]);
  assign t[35] = t[3] ? t[38] : t[37];
  assign t[36] = ~(t[6] & t[62]);
  assign t[37] = ~(t[63]);
  assign t[38] = ~(t[54] & t[39]);
  assign t[39] = x[18] ? x[34] : t[40];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[41] | t[42]);
  assign t[41] = ~(t[30] | t[31]);
  assign t[42] = ~(t[17] | t[43]);
  assign t[43] = ~(t[56] ^ t[58]);
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[64]);
  assign t[47] = ~(t[65]);
  assign t[48] = ~(t[54] & t[49]);
  assign t[49] = x[18] ? x[37] : t[50];
  assign t[4] = ~(t[53]);
  assign t[50] = ~(t[51] ^ t[43]);
  assign t[51] = ~(t[17] | t[57]);
  assign t[52] = (t[66]);
  assign t[53] = (t[67]);
  assign t[54] = (t[68]);
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[54] & t[8]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = t[80] ^ x[5];
  assign t[67] = t[81] ^ x[11];
  assign t[68] = t[82] ^ x[14];
  assign t[69] = t[83] ^ x[17];
  assign t[6] = ~(t[54] | t[7]);
  assign t[70] = t[84] ^ x[25];
  assign t[71] = t[85] ^ x[26];
  assign t[72] = t[86] ^ x[27];
  assign t[73] = t[87] ^ x[28];
  assign t[74] = t[88] ^ x[29];
  assign t[75] = t[89] ^ x[30];
  assign t[76] = t[90] ^ x[32];
  assign t[77] = t[91] ^ x[33];
  assign t[78] = t[92] ^ x[35];
  assign t[79] = t[93] ^ x[36];
  assign t[7] = ~(t[55]);
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[102] & t[104]);
  assign t[86] = (~t[102] & t[105]);
  assign t[87] = (~t[102] & t[106]);
  assign t[88] = (~t[94] & t[107]);
  assign t[89] = (~t[96] & t[108]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[90] = (~t[94] & t[109]);
  assign t[91] = (~t[96] & t[110]);
  assign t[92] = (~t[94] & t[111]);
  assign t[93] = (~t[96] & t[112]);
  assign t[94] = t[113] ^ x[4];
  assign t[95] = t[114] ^ x[5];
  assign t[96] = t[115] ^ x[10];
  assign t[97] = t[116] ^ x[11];
  assign t[98] = t[117] ^ x[13];
  assign t[99] = t[118] ^ x[14];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0] & ~t[20] & ~t[34] & ~t[44]) | (~t[0] & t[20] & ~t[34] & ~t[44]) | (~t[0] & ~t[20] & t[34] & ~t[44]) | (~t[0] & ~t[20] & ~t[34] & t[44]) | (t[0] & t[20] & t[34] & ~t[44]) | (t[0] & t[20] & ~t[34] & t[44]) | (t[0] & ~t[20] & t[34] & t[44]) | (~t[0] & t[20] & t[34] & t[44]);
endmodule

module R2ind311(x, y);
 input [28:0] x;
 output y;

 wire [62:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[17]);
  assign t[11] = ~(t[18] ^ t[19]);
  assign t[12] = ~(t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = t[29] ^ x[5];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = t[31] ^ x[14];
  assign t[24] = t[32] ^ x[17];
  assign t[25] = t[33] ^ x[25];
  assign t[26] = t[34] ^ x[26];
  assign t[27] = t[35] ^ x[27];
  assign t[28] = t[36] ^ x[28];
  assign t[29] = (~t[37] & t[38]);
  assign t[2] = ~(t[6] & t[13]);
  assign t[30] = (~t[39] & t[40]);
  assign t[31] = (~t[41] & t[42]);
  assign t[32] = (~t[43] & t[44]);
  assign t[33] = (~t[45] & t[46]);
  assign t[34] = (~t[45] & t[47]);
  assign t[35] = (~t[45] & t[48]);
  assign t[36] = (~t[45] & t[49]);
  assign t[37] = t[50] ^ x[4];
  assign t[38] = t[51] ^ x[5];
  assign t[39] = t[52] ^ x[10];
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] ^ x[11];
  assign t[41] = t[54] ^ x[13];
  assign t[42] = t[55] ^ x[14];
  assign t[43] = t[56] ^ x[16];
  assign t[44] = t[57] ^ x[17];
  assign t[45] = t[58] ^ x[24];
  assign t[46] = t[59] ^ x[25];
  assign t[47] = t[60] ^ x[26];
  assign t[48] = t[61] ^ x[27];
  assign t[49] = t[62] ^ x[28];
  assign t[4] = ~(t[14]);
  assign t[50] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[51] = (x[3]);
  assign t[52] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[53] = (x[9]);
  assign t[54] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[12]);
  assign t[56] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[15]);
  assign t[58] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[59] = (x[21]);
  assign t[5] = ~(t[15] & t[8]);
  assign t[60] = (x[23]);
  assign t[61] = (x[20]);
  assign t[62] = (x[22]);
  assign t[6] = ~(t[15] | t[7]);
  assign t[7] = ~(t[16]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = ~(t[10] ^ t[11]);
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [28:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[14]);
  assign t[13] = t[24] ? t[17] : t[25];
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[24] ^ t[27]);
  assign t[16] = ~(t[24] | t[27]);
  assign t[17] = ~(t[25] & t[18]);
  assign t[18] = ~(t[19] & t[14]);
  assign t[19] = ~(t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[5];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[14];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[25];
  assign t[33] = t[41] ^ x[26];
  assign t[34] = t[42] ^ x[27];
  assign t[35] = t[43] ^ x[28];
  assign t[36] = (~t[44] & t[45]);
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[52] & t[54]);
  assign t[42] = (~t[52] & t[55]);
  assign t[43] = (~t[52] & t[56]);
  assign t[44] = t[57] ^ x[4];
  assign t[45] = t[58] ^ x[5];
  assign t[46] = t[59] ^ x[10];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[13];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~(t[21]);
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[17];
  assign t[52] = t[65] ^ x[24];
  assign t[53] = t[66] ^ x[25];
  assign t[54] = t[67] ^ x[26];
  assign t[55] = t[68] ^ x[27];
  assign t[56] = t[69] ^ x[28];
  assign t[57] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[58] = (x[2]);
  assign t[59] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[8]);
  assign t[61] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[12]);
  assign t[63] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[15]);
  assign t[65] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[66] = (x[23]);
  assign t[67] = (x[21]);
  assign t[68] = (x[22]);
  assign t[69] = (x[20]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = ~(t[10] | t[11]);
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [28:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[28] | t[16]);
  assign t[13] = ~(t[29] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = t[30] ? t[13] : t[29];
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[22] & t[19]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[29]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[6] & t[24]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[11];
  assign t[34] = t[42] ^ x[14];
  assign t[35] = t[43] ^ x[17];
  assign t[36] = t[44] ^ x[25];
  assign t[37] = t[45] ^ x[26];
  assign t[38] = t[46] ^ x[27];
  assign t[39] = t[47] ^ x[28];
  assign t[3] = ~(t[7]);
  assign t[40] = (~t[48] & t[49]);
  assign t[41] = (~t[50] & t[51]);
  assign t[42] = (~t[52] & t[53]);
  assign t[43] = (~t[54] & t[55]);
  assign t[44] = (~t[56] & t[57]);
  assign t[45] = (~t[56] & t[58]);
  assign t[46] = (~t[56] & t[59]);
  assign t[47] = (~t[56] & t[60]);
  assign t[48] = t[61] ^ x[4];
  assign t[49] = t[62] ^ x[5];
  assign t[4] = ~(t[25]);
  assign t[50] = t[63] ^ x[10];
  assign t[51] = t[64] ^ x[11];
  assign t[52] = t[65] ^ x[13];
  assign t[53] = t[66] ^ x[14];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[17];
  assign t[56] = t[69] ^ x[24];
  assign t[57] = t[70] ^ x[25];
  assign t[58] = t[71] ^ x[26];
  assign t[59] = t[72] ^ x[27];
  assign t[5] = ~(t[26] & t[8]);
  assign t[60] = t[73] ^ x[28];
  assign t[61] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[62] = (x[1]);
  assign t[63] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[64] = (x[7]);
  assign t[65] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[12]);
  assign t[67] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[15]);
  assign t[69] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[6] = ~(t[26] | t[7]);
  assign t[70] = (x[22]);
  assign t[71] = (x[21]);
  assign t[72] = (x[23]);
  assign t[73] = (x[20]);
  assign t[7] = ~(t[27]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [28:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[24] ? t[13] : t[12];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[25] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[24] | t[26]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[19] & t[17]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[19] & t[15]);
  assign t[19] = ~(t[26]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[5];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[14];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[25];
  assign t[33] = t[41] ^ x[26];
  assign t[34] = t[42] ^ x[27];
  assign t[35] = t[43] ^ x[28];
  assign t[36] = (~t[44] & t[45]);
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[52] & t[54]);
  assign t[42] = (~t[52] & t[55]);
  assign t[43] = (~t[52] & t[56]);
  assign t[44] = t[57] ^ x[4];
  assign t[45] = t[58] ^ x[5];
  assign t[46] = t[59] ^ x[10];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[13];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~(t[21]);
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[17];
  assign t[52] = t[65] ^ x[24];
  assign t[53] = t[66] ^ x[25];
  assign t[54] = t[67] ^ x[26];
  assign t[55] = t[68] ^ x[27];
  assign t[56] = t[69] ^ x[28];
  assign t[57] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[58] = (x[0]);
  assign t[59] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[6]);
  assign t[61] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[12]);
  assign t[63] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[15]);
  assign t[65] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[66] = (x[23]);
  assign t[67] = (x[21]);
  assign t[68] = (x[20]);
  assign t[69] = (x[22]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[18] ? x[19] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [37:0] x;
 output y;

 wire [102:0] t;
  assign t[0] = t[1] ? t[14] : t[2];
  assign t[100] = (x[8]);
  assign t[101] = (x[26]);
  assign t[102] = (x[7]);
  assign t[10] = t[1] ? t[24] : t[11];
  assign t[11] = t[25] ^ t[26];
  assign t[12] = t[1] ? t[27] : t[13];
  assign t[13] = t[14] ^ t[28];
  assign t[14] = (t[29]);
  assign t[15] = (t[30]);
  assign t[16] = (t[31]);
  assign t[17] = (t[32]);
  assign t[18] = (t[33]);
  assign t[19] = (t[34]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[35]);
  assign t[21] = (t[36]);
  assign t[22] = (t[37]);
  assign t[23] = (t[38]);
  assign t[24] = (t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = t[44] ^ x[5];
  assign t[2] = t[15] ^ t[16];
  assign t[30] = t[45] ^ x[6];
  assign t[31] = t[46] ^ x[12];
  assign t[32] = t[47] ^ x[15];
  assign t[33] = t[48] ^ x[18];
  assign t[34] = t[49] ^ x[21];
  assign t[35] = t[50] ^ x[24];
  assign t[36] = t[51] ^ x[30];
  assign t[37] = t[52] ^ x[31];
  assign t[38] = t[53] ^ x[32];
  assign t[39] = t[54] ^ x[33];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[55] ^ x[34];
  assign t[41] = t[56] ^ x[35];
  assign t[42] = t[57] ^ x[36];
  assign t[43] = t[58] ^ x[37];
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[59] & t[61]);
  assign t[46] = (~t[62] & t[63]);
  assign t[47] = (~t[64] & t[65]);
  assign t[48] = (~t[66] & t[67]);
  assign t[49] = (~t[68] & t[69]);
  assign t[4] = ~(t[17] & t[7]);
  assign t[50] = (~t[70] & t[71]);
  assign t[51] = (~t[72] & t[73]);
  assign t[52] = (~t[59] & t[74]);
  assign t[53] = (~t[62] & t[75]);
  assign t[54] = (~t[72] & t[76]);
  assign t[55] = (~t[59] & t[77]);
  assign t[56] = (~t[62] & t[78]);
  assign t[57] = (~t[72] & t[79]);
  assign t[58] = (~t[62] & t[80]);
  assign t[59] = t[81] ^ x[4];
  assign t[5] = ~(t[18]);
  assign t[60] = t[82] ^ x[5];
  assign t[61] = t[83] ^ x[6];
  assign t[62] = t[84] ^ x[11];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[15];
  assign t[66] = t[88] ^ x[17];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[20];
  assign t[69] = t[91] ^ x[21];
  assign t[6] = ~(t[19]);
  assign t[70] = t[92] ^ x[23];
  assign t[71] = t[93] ^ x[24];
  assign t[72] = t[94] ^ x[29];
  assign t[73] = t[95] ^ x[30];
  assign t[74] = t[96] ^ x[31];
  assign t[75] = t[97] ^ x[32];
  assign t[76] = t[98] ^ x[33];
  assign t[77] = t[99] ^ x[34];
  assign t[78] = t[100] ^ x[35];
  assign t[79] = t[101] ^ x[36];
  assign t[7] = ~(t[20]);
  assign t[80] = t[102] ^ x[37];
  assign t[81] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[82] = (x[0]);
  assign t[83] = (x[3]);
  assign t[84] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[85] = (x[10]);
  assign t[86] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[13]);
  assign t[88] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[16]);
  assign t[8] = t[1] ? t[21] : t[9];
  assign t[90] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[19]);
  assign t[92] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[22]);
  assign t[94] = (x[25] & ~x[26] & ~x[27] & ~x[28]) | (~x[25] & x[26] & ~x[27] & ~x[28]) | (~x[25] & ~x[26] & x[27] & ~x[28]) | (~x[25] & ~x[26] & ~x[27] & x[28]) | (x[25] & x[26] & x[27] & ~x[28]) | (x[25] & x[26] & ~x[27] & x[28]) | (x[25] & ~x[26] & x[27] & x[28]) | (~x[25] & x[26] & x[27] & x[28]);
  assign t[95] = (x[28]);
  assign t[96] = (x[2]);
  assign t[97] = (x[9]);
  assign t[98] = (x[27]);
  assign t[99] = (x[1]);
  assign t[9] = t[22] ^ t[23];
  assign y = (t[0] & ~t[8] & ~t[10] & ~t[12]) | (~t[0] & t[8] & ~t[10] & ~t[12]) | (~t[0] & ~t[8] & t[10] & ~t[12]) | (~t[0] & ~t[8] & ~t[10] & t[12]) | (t[0] & t[8] & t[10] & ~t[12]) | (t[0] & t[8] & ~t[10] & t[12]) | (t[0] & ~t[8] & t[10] & t[12]) | (~t[0] & t[8] & t[10] & t[12]);
endmodule

module R2ind316(x, y);
 input [29:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[5];
  assign t[16] = t[23] ^ x[11];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[20];
  assign t[19] = t[26] ^ x[23];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[29];
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = (~t[35] & t[36]);
  assign t[26] = (~t[37] & t[38]);
  assign t[27] = (~t[39] & t[40]);
  assign t[28] = (~t[41] & t[42]);
  assign t[29] = t[43] ^ x[4];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[5];
  assign t[31] = t[45] ^ x[10];
  assign t[32] = t[46] ^ x[11];
  assign t[33] = t[47] ^ x[16];
  assign t[34] = t[48] ^ x[17];
  assign t[35] = t[49] ^ x[19];
  assign t[36] = t[50] ^ x[20];
  assign t[37] = t[51] ^ x[22];
  assign t[38] = t[52] ^ x[23];
  assign t[39] = t[53] ^ x[25];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[26];
  assign t[41] = t[55] ^ x[28];
  assign t[42] = t[56] ^ x[29];
  assign t[43] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[44] = (x[1]);
  assign t[45] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[46] = (x[6]);
  assign t[47] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[48] = (x[12]);
  assign t[49] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[18]);
  assign t[51] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[21]);
  assign t[53] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[24]);
  assign t[55] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[27]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [29:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[5];
  assign t[16] = t[23] ^ x[11];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[20];
  assign t[19] = t[26] ^ x[23];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[29];
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = (~t[35] & t[36]);
  assign t[26] = (~t[37] & t[38]);
  assign t[27] = (~t[39] & t[40]);
  assign t[28] = (~t[41] & t[42]);
  assign t[29] = t[43] ^ x[4];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[5];
  assign t[31] = t[45] ^ x[10];
  assign t[32] = t[46] ^ x[11];
  assign t[33] = t[47] ^ x[16];
  assign t[34] = t[48] ^ x[17];
  assign t[35] = t[49] ^ x[19];
  assign t[36] = t[50] ^ x[20];
  assign t[37] = t[51] ^ x[22];
  assign t[38] = t[52] ^ x[23];
  assign t[39] = t[53] ^ x[25];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[26];
  assign t[41] = t[55] ^ x[28];
  assign t[42] = t[56] ^ x[29];
  assign t[43] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[44] = (x[2]);
  assign t[45] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[46] = (x[7]);
  assign t[47] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[48] = (x[13]);
  assign t[49] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[18]);
  assign t[51] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[21]);
  assign t[53] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[24]);
  assign t[55] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[27]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [29:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[5];
  assign t[16] = t[23] ^ x[11];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[20];
  assign t[19] = t[26] ^ x[23];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[29];
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[31] & t[32]);
  assign t[24] = (~t[33] & t[34]);
  assign t[25] = (~t[35] & t[36]);
  assign t[26] = (~t[37] & t[38]);
  assign t[27] = (~t[39] & t[40]);
  assign t[28] = (~t[41] & t[42]);
  assign t[29] = t[43] ^ x[4];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[5];
  assign t[31] = t[45] ^ x[10];
  assign t[32] = t[46] ^ x[11];
  assign t[33] = t[47] ^ x[16];
  assign t[34] = t[48] ^ x[17];
  assign t[35] = t[49] ^ x[19];
  assign t[36] = t[50] ^ x[20];
  assign t[37] = t[51] ^ x[22];
  assign t[38] = t[52] ^ x[23];
  assign t[39] = t[53] ^ x[25];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[26];
  assign t[41] = t[55] ^ x[28];
  assign t[42] = t[56] ^ x[29];
  assign t[43] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[44] = (x[3]);
  assign t[45] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[46] = (x[8]);
  assign t[47] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[48] = (x[14]);
  assign t[49] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[18]);
  assign t[51] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[21]);
  assign t[53] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[24]);
  assign t[55] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[27]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [24:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[5];
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[12];
  assign t[18] = t[25] ^ x[15];
  assign t[19] = t[26] ^ x[18];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[21];
  assign t[21] = t[28] ^ x[24];
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[29] & t[31]);
  assign t[24] = (~t[32] & t[33]);
  assign t[25] = (~t[34] & t[35]);
  assign t[26] = (~t[36] & t[37]);
  assign t[27] = (~t[38] & t[39]);
  assign t[28] = (~t[40] & t[41]);
  assign t[29] = t[42] ^ x[4];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[43] ^ x[5];
  assign t[31] = t[44] ^ x[6];
  assign t[32] = t[45] ^ x[11];
  assign t[33] = t[46] ^ x[12];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[15];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[18];
  assign t[38] = t[51] ^ x[20];
  assign t[39] = t[52] ^ x[21];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[24];
  assign t[42] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[43] = (x[0]);
  assign t[44] = (x[3]);
  assign t[45] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[46] = (x[10]);
  assign t[47] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[48] = (x[13]);
  assign t[49] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[16]);
  assign t[51] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[19]);
  assign t[53] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[22]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [558:0] x;
 output [319:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[33]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[33]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[8], x[7], x[6], x[17], x[16], x[15], x[33]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[8], x[7], x[6], x[17], x[16], x[15], x[33]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[36], x[35], x[34], x[42], x[41], x[40], x[39], x[38], x[37], x[33], x[45], x[44], x[43]}), .y(y[30]));
  R2ind31 R2ind31_inst(.y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[36], x[35], x[34], x[42], x[41], x[40], x[39], x[38], x[37], x[33], x[45], x[44], x[43]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[33], x[36], x[35], x[34], x[42], x[41], x[40]}), .y(y[35]));
  R2ind36 R2ind36_inst(.y(y[36]));
  R2ind37 R2ind37_inst(.y(y[37]));
  R2ind38 R2ind38_inst(.y(y[38]));
  R2ind39 R2ind39_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[33], x[36], x[35], x[34], x[42], x[41], x[40]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33], x[48], x[47], x[46], x[36], x[35], x[34]}), .y(y[40]));
  R2ind41 R2ind41_inst(.y(y[41]));
  R2ind42 R2ind42_inst(.y(y[42]));
  R2ind43 R2ind43_inst(.y(y[43]));
  R2ind44 R2ind44_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33], x[48], x[47], x[46], x[36], x[35], x[34]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33], x[48], x[47], x[46]}), .y(y[45]));
  R2ind46 R2ind46_inst(.y(y[46]));
  R2ind47 R2ind47_inst(.y(y[47]));
  R2ind48 R2ind48_inst(.y(y[48]));
  R2ind49 R2ind49_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[33], x[48], x[47], x[46]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[36], x[35], x[34], x[42], x[41], x[40], x[33], x[39], x[38], x[37]}), .y(y[50]));
  R2ind51 R2ind51_inst(.y(y[51]));
  R2ind52 R2ind52_inst(.y(y[52]));
  R2ind53 R2ind53_inst(.y(y[53]));
  R2ind54 R2ind54_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[48], x[47], x[46], x[36], x[35], x[34], x[42], x[41], x[40], x[33], x[39], x[38], x[37]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[32], x[31], x[30], x[51], x[50], x[49], x[23], x[22], x[21]}), .y(y[55]));
  R2ind56 R2ind56_inst(.y(y[56]));
  R2ind57 R2ind57_inst(.y(y[57]));
  R2ind58 R2ind58_inst(.y(y[58]));
  R2ind59 R2ind59_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[32], x[31], x[30], x[51], x[50], x[49], x[23], x[22], x[21]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[32], x[31], x[30], x[23], x[22], x[21], x[51], x[50], x[49], x[26], x[25], x[24]}), .y(y[60]));
  R2ind61 R2ind61_inst(.y(y[61]));
  R2ind62 R2ind62_inst(.y(y[62]));
  R2ind63 R2ind63_inst(.y(y[63]));
  R2ind64 R2ind64_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[32], x[31], x[30], x[23], x[22], x[21], x[51], x[50], x[49], x[26], x[25], x[24]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[51], x[50], x[49], x[32], x[31], x[30]}), .y(y[65]));
  R2ind66 R2ind66_inst(.y(y[66]));
  R2ind67 R2ind67_inst(.y(y[67]));
  R2ind68 R2ind68_inst(.y(y[68]));
  R2ind69 R2ind69_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[51], x[50], x[49], x[32], x[31], x[30]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[51], x[50], x[49]}), .y(y[70]));
  R2ind71 R2ind71_inst(.y(y[71]));
  R2ind72 R2ind72_inst(.y(y[72]));
  R2ind73 R2ind73_inst(.y(y[73]));
  R2ind74 R2ind74_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[8], x[7], x[6], x[29], x[28], x[27], x[51], x[50], x[49]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[17], x[16], x[15], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9]}), .y(y[75]));
  R2ind76 R2ind76_inst(.y(y[76]));
  R2ind77 R2ind77_inst(.y(y[77]));
  R2ind78 R2ind78_inst(.y(y[78]));
  R2ind79 R2ind79_inst(.x({x[17], x[16], x[15], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[33]}), .y(y[80]));
  R2ind81 R2ind81_inst(.y(y[81]));
  R2ind82 R2ind82_inst(.y(y[82]));
  R2ind83 R2ind83_inst(.y(y[83]));
  R2ind84 R2ind84_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[33]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[51], x[50], x[49], x[8], x[7], x[6]}), .y(y[85]));
  R2ind86 R2ind86_inst(.y(y[86]));
  R2ind87 R2ind87_inst(.y(y[87]));
  R2ind88 R2ind88_inst(.y(y[88]));
  R2ind89 R2ind89_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[20], x[19], x[18], x[51], x[50], x[49], x[8], x[7], x[6]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[51], x[50], x[49]}), .y(y[90]));
  R2ind91 R2ind91_inst(.y(y[91]));
  R2ind92 R2ind92_inst(.y(y[92]));
  R2ind93 R2ind93_inst(.y(y[93]));
  R2ind94 R2ind94_inst(.x({x[51], x[50], x[49]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[51], x[50], x[49]}), .y(y[95]));
  R2ind96 R2ind96_inst(.y(y[96]));
  R2ind97 R2ind97_inst(.y(y[97]));
  R2ind98 R2ind98_inst(.y(y[98]));
  R2ind99 R2ind99_inst(.x({x[51], x[50], x[49]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[54], x[53], x[52]}), .y(y[100]));
  R2ind101 R2ind101_inst(.y(y[101]));
  R2ind102 R2ind102_inst(.y(y[102]));
  R2ind103 R2ind103_inst(.y(y[103]));
  R2ind104 R2ind104_inst(.x({x[54], x[53], x[52]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[54], x[53], x[52]}), .y(y[105]));
  R2ind106 R2ind106_inst(.y(y[106]));
  R2ind107 R2ind107_inst(.y(y[107]));
  R2ind108 R2ind108_inst(.y(y[108]));
  R2ind109 R2ind109_inst(.x({x[54], x[53], x[52]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[57], x[56], x[55]}), .y(y[110]));
  R2ind111 R2ind111_inst(.y(y[111]));
  R2ind112 R2ind112_inst(.y(y[112]));
  R2ind113 R2ind113_inst(.y(y[113]));
  R2ind114 R2ind114_inst(.x({x[57], x[56], x[55]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[60], x[59], x[58]}), .y(y[115]));
  R2ind116 R2ind116_inst(.y(y[116]));
  R2ind117 R2ind117_inst(.y(y[117]));
  R2ind118 R2ind118_inst(.y(y[118]));
  R2ind119 R2ind119_inst(.x({x[60], x[59], x[58]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[60], x[59], x[58]}), .y(y[120]));
  R2ind121 R2ind121_inst(.y(y[121]));
  R2ind122 R2ind122_inst(.y(y[122]));
  R2ind123 R2ind123_inst(.y(y[123]));
  R2ind124 R2ind124_inst(.x({x[60], x[59], x[58]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[63], x[62], x[61]}), .y(y[125]));
  R2ind126 R2ind126_inst(.y(y[126]));
  R2ind127 R2ind127_inst(.y(y[127]));
  R2ind128 R2ind128_inst(.y(y[128]));
  R2ind129 R2ind129_inst(.x({x[63], x[62], x[61]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[63], x[62], x[61]}), .y(y[130]));
  R2ind131 R2ind131_inst(.y(y[131]));
  R2ind132 R2ind132_inst(.y(y[132]));
  R2ind133 R2ind133_inst(.y(y[133]));
  R2ind134 R2ind134_inst(.x({x[63], x[62], x[61]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[33], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[8], x[7], x[6], x[51], x[50], x[49], x[69], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[91], x[90], x[88], x[33], x[89], x[87], x[86], x[85], x[84], x[83], x[121], x[81], x[80], x[79], x[78], x[77], x[120], x[75], x[74], x[73], x[72], x[71], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[8], x[7], x[6], x[51], x[50], x[49], x[112], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[90], x[89], x[88], x[91], x[87], x[86], x[85], x[84], x[83], x[33], x[111], x[81], x[80], x[79], x[78], x[77], x[110], x[75], x[74], x[73], x[72], x[71], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[8], x[7], x[6], x[51], x[50], x[49], x[102], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[90], x[91], x[88], x[89], x[87], x[86], x[85], x[84], x[83], x[33], x[101], x[81], x[80], x[79], x[78], x[77], x[100], x[75], x[74], x[73], x[72], x[71], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[8], x[7], x[6], x[51], x[50], x[49], x[92], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[91], x[33], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[8], x[7], x[6], x[51], x[50], x[49], x[69], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[98], x[69], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[92], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[102], x[33], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[57], x[56], x[55], x[51], x[50], x[49], x[122], x[97], x[96], x[95], x[94], x[93], x[112], x[68], x[67], x[66], x[65], x[64]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[33], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[57], x[56], x[55], x[51], x[50], x[49], x[98], x[97], x[96], x[95], x[94], x[93], x[69], x[68], x[67], x[66], x[65], x[64]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[57], x[56], x[55], x[51], x[50], x[49], x[138], x[97], x[96], x[95], x[94], x[93], x[92], x[68], x[67], x[66], x[65], x[64]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[33], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[57], x[56], x[55], x[51], x[50], x[49], x[130], x[97], x[96], x[95], x[94], x[93], x[102], x[68], x[67], x[66], x[65], x[64]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[33], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[57], x[56], x[55], x[51], x[50], x[49], x[122], x[97], x[96], x[95], x[94], x[93], x[112], x[68], x[67], x[66], x[65], x[64]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[108], x[98], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[138], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[130], x[33], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[57], x[56], x[55], x[156], x[155], x[154], x[153], x[107], x[106], x[105], x[104], x[103], x[122], x[97], x[96], x[95], x[94], x[93]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[33], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55], x[156], x[155], x[154], x[108], x[107], x[106], x[105], x[104], x[103], x[98], x[97], x[96], x[95], x[94], x[93]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[33], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55], x[156], x[155], x[154], x[172], x[107], x[106], x[105], x[104], x[103], x[138], x[97], x[96], x[95], x[94], x[93]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[33], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55], x[156], x[155], x[154], x[164], x[107], x[106], x[105], x[104], x[103], x[130], x[97], x[96], x[95], x[94], x[93]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[33], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[57], x[56], x[55], x[156], x[155], x[154], x[153], x[107], x[106], x[105], x[104], x[103], x[122], x[97], x[96], x[95], x[94], x[93]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[118], x[108], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[172], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[164], x[33], x[188], x[82], x[81], x[80], x[79], x[78], x[77], x[57], x[56], x[55], x[156], x[155], x[154], x[187], x[117], x[116], x[115], x[114], x[113], x[153], x[107], x[106], x[105], x[104], x[103]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[33], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[57], x[56], x[55], x[156], x[155], x[154], x[118], x[117], x[116], x[115], x[114], x[113], x[108], x[107], x[106], x[105], x[104], x[103]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[33], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[57], x[56], x[55], x[156], x[155], x[154], x[197], x[117], x[116], x[115], x[114], x[113], x[172], x[107], x[106], x[105], x[104], x[103]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[33], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[57], x[56], x[55], x[156], x[155], x[154], x[189], x[117], x[116], x[115], x[114], x[113], x[164], x[107], x[106], x[105], x[104], x[103]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[33], x[188], x[82], x[81], x[80], x[79], x[78], x[77], x[57], x[56], x[55], x[156], x[155], x[154], x[187], x[117], x[116], x[115], x[114], x[113], x[153], x[107], x[106], x[105], x[104], x[103]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[218], x[92], x[68], x[67], x[66], x[65], x[64], x[151], x[118], x[217], x[138], x[97], x[96], x[95], x[94], x[93], x[216], x[215], x[172], x[107], x[106], x[105], x[104], x[103], x[214], x[189], x[33], x[213], x[197], x[156], x[155], x[154], x[212], x[150], x[149], x[148], x[147], x[146], x[187], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[33], x[218], x[92], x[68], x[67], x[66], x[65], x[64], x[156], x[155], x[154], x[151], x[150], x[149], x[148], x[147], x[146], x[118], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[33], x[217], x[138], x[97], x[96], x[95], x[94], x[93], x[156], x[155], x[154], x[216], x[150], x[149], x[148], x[147], x[146], x[197], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[33], x[215], x[172], x[107], x[106], x[105], x[104], x[103], x[156], x[155], x[154], x[214], x[150], x[149], x[148], x[147], x[146], x[189], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[33], x[213], x[197], x[156], x[155], x[154], x[212], x[150], x[149], x[148], x[147], x[146], x[187], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[227], x[144], x[151], x[226], x[225], x[216], x[224], x[223], x[135], x[134], x[133], x[132], x[131], x[222], x[214], x[33], x[221], x[220], x[127], x[126], x[125], x[124], x[123], x[57], x[56], x[55], x[156], x[155], x[154], x[219], x[143], x[142], x[141], x[140], x[139], x[212], x[150], x[149], x[148], x[147], x[146]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[33], x[227], x[216], x[57], x[56], x[55], x[156], x[155], x[154], x[144], x[143], x[142], x[141], x[140], x[139], x[151], x[150], x[149], x[148], x[147], x[146]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[33], x[226], x[57], x[56], x[55], x[156], x[155], x[154], x[225], x[143], x[142], x[141], x[140], x[139], x[216], x[150], x[149], x[148], x[147], x[146]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[33], x[224], x[223], x[135], x[134], x[133], x[132], x[131], x[57], x[56], x[55], x[156], x[155], x[154], x[222], x[143], x[142], x[141], x[140], x[139], x[214], x[150], x[149], x[148], x[147], x[146]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[33], x[221], x[220], x[127], x[126], x[125], x[124], x[123], x[57], x[56], x[55], x[156], x[155], x[154], x[219], x[143], x[142], x[141], x[140], x[139], x[212], x[150], x[149], x[148], x[147], x[146]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[237], x[236], x[184], x[183], x[182], x[181], x[180], x[136], x[144], x[235], x[234], x[177], x[176], x[175], x[174], x[173], x[223], x[225], x[233], x[232], x[169], x[168], x[167], x[166], x[165], x[231], x[222], x[33], x[230], x[229], x[161], x[160], x[159], x[158], x[157], x[57], x[56], x[55], x[156], x[155], x[154], x[228], x[135], x[134], x[133], x[132], x[131], x[219], x[143], x[142], x[141], x[140], x[139]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[33], x[237], x[236], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55], x[156], x[155], x[154], x[136], x[135], x[134], x[133], x[132], x[131], x[144], x[143], x[142], x[141], x[140], x[139]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[33], x[235], x[234], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55], x[156], x[155], x[154], x[223], x[135], x[134], x[133], x[132], x[131], x[225], x[143], x[142], x[141], x[140], x[139]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[33], x[233], x[232], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55], x[156], x[155], x[154], x[231], x[135], x[134], x[133], x[132], x[131], x[222], x[143], x[142], x[141], x[140], x[139]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[33], x[230], x[229], x[161], x[160], x[159], x[158], x[157], x[57], x[56], x[55], x[156], x[155], x[154], x[228], x[135], x[134], x[133], x[132], x[131], x[219], x[143], x[142], x[141], x[140], x[139]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[246], x[245], x[209], x[208], x[207], x[206], x[205], x[128], x[136], x[244], x[243], x[202], x[201], x[200], x[199], x[198], x[220], x[223], x[242], x[241], x[194], x[193], x[192], x[191], x[190], x[240], x[231], x[33], x[239], x[101], x[81], x[80], x[79], x[78], x[77], x[57], x[56], x[55], x[156], x[155], x[154], x[238], x[127], x[126], x[125], x[124], x[123], x[228], x[135], x[134], x[133], x[132], x[131]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[33], x[246], x[245], x[209], x[208], x[207], x[206], x[205], x[57], x[56], x[55], x[156], x[155], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[136], x[135], x[134], x[133], x[132], x[131]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[33], x[244], x[243], x[202], x[201], x[200], x[199], x[198], x[57], x[56], x[55], x[156], x[155], x[154], x[220], x[127], x[126], x[125], x[124], x[123], x[223], x[135], x[134], x[133], x[132], x[131]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[33], x[242], x[241], x[194], x[193], x[192], x[191], x[190], x[57], x[56], x[55], x[156], x[155], x[154], x[240], x[127], x[126], x[125], x[124], x[123], x[231], x[135], x[134], x[133], x[132], x[131]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[33], x[239], x[101], x[81], x[80], x[79], x[78], x[77], x[57], x[56], x[55], x[156], x[155], x[154], x[238], x[127], x[126], x[125], x[124], x[123], x[228], x[135], x[134], x[133], x[132], x[131]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[252], x[102], x[68], x[67], x[66], x[65], x[64], x[185], x[128], x[251], x[130], x[97], x[96], x[95], x[94], x[93], x[236], x[220], x[250], x[164], x[107], x[106], x[105], x[104], x[103], x[249], x[240], x[33], x[248], x[189], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55], x[156], x[155], x[154], x[247], x[184], x[183], x[182], x[181], x[180], x[238], x[127], x[126], x[125], x[124], x[123]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[33], x[252], x[102], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55], x[156], x[155], x[154], x[185], x[184], x[183], x[182], x[181], x[180], x[128], x[127], x[126], x[125], x[124], x[123]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[33], x[251], x[130], x[97], x[96], x[95], x[94], x[93], x[57], x[56], x[55], x[156], x[155], x[154], x[236], x[184], x[183], x[182], x[181], x[180], x[220], x[127], x[126], x[125], x[124], x[123]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[33], x[250], x[164], x[107], x[106], x[105], x[104], x[103], x[57], x[56], x[55], x[156], x[155], x[154], x[249], x[184], x[183], x[182], x[181], x[180], x[240], x[127], x[126], x[125], x[124], x[123]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[33], x[248], x[189], x[117], x[116], x[115], x[114], x[113], x[57], x[56], x[55], x[156], x[155], x[154], x[247], x[184], x[183], x[182], x[181], x[180], x[238], x[127], x[126], x[125], x[124], x[123]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[261], x[214], x[150], x[149], x[148], x[147], x[146], x[178], x[185], x[260], x[222], x[143], x[142], x[141], x[140], x[139], x[234], x[236], x[259], x[231], x[135], x[134], x[133], x[132], x[131], x[258], x[249], x[257], x[240], x[127], x[126], x[125], x[124], x[123], x[33], x[256], x[255], x[254], x[253], x[177], x[176], x[175], x[174], x[173], x[247], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[33], x[261], x[214], x[150], x[149], x[148], x[147], x[146], x[256], x[255], x[254], x[178], x[177], x[176], x[175], x[174], x[173], x[185], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[33], x[260], x[222], x[143], x[142], x[141], x[140], x[139], x[256], x[255], x[254], x[234], x[177], x[176], x[175], x[174], x[173], x[236], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[33], x[259], x[231], x[135], x[134], x[133], x[132], x[131], x[256], x[255], x[254], x[258], x[177], x[176], x[175], x[174], x[173], x[249], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[257], x[240], x[127], x[126], x[125], x[124], x[123], x[33], x[256], x[255], x[254], x[253], x[177], x[176], x[175], x[174], x[173], x[247], x[184], x[183], x[182], x[181], x[180], x[57], x[56], x[55]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[288], x[287], x[76], x[286], x[285], x[284], x[100], x[283], x[282], x[281], x[110], x[280], x[279], x[278], x[277], x[276], x[275], x[274], x[33], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[120], x[75], x[74], x[73], x[72], x[71], x[264], x[263], x[262]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[288], x[270], x[33], x[273], x[272], x[271], x[287], x[269], x[268], x[267], x[266], x[265], x[76], x[75], x[74], x[73], x[72], x[71], x[264], x[263], x[262]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[286], x[285], x[278], x[277], x[276], x[275], x[274], x[33], x[273], x[272], x[271], x[284], x[269], x[268], x[267], x[266], x[265], x[100], x[75], x[74], x[73], x[72], x[71], x[264], x[263], x[262]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[283], x[282], x[278], x[277], x[276], x[275], x[274], x[33], x[273], x[272], x[271], x[281], x[269], x[268], x[267], x[266], x[265], x[110], x[75], x[74], x[73], x[72], x[71], x[264], x[263], x[262]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[280], x[279], x[278], x[277], x[276], x[275], x[274], x[33], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[120], x[75], x[74], x[73], x[72], x[71], x[264], x[263], x[262]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[304], x[285], x[287], x[303], x[302], x[282], x[284], x[301], x[300], x[279], x[281], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[33], x[292], x[291], x[290], x[289], x[278], x[277], x[276], x[275], x[274], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[304], x[289], x[33], x[292], x[291], x[290], x[285], x[278], x[277], x[276], x[275], x[274], x[287], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[303], x[302], x[297], x[296], x[295], x[294], x[293], x[33], x[292], x[291], x[290], x[282], x[278], x[277], x[276], x[275], x[274], x[284], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[301], x[300], x[297], x[296], x[295], x[294], x[293], x[33], x[292], x[291], x[290], x[279], x[278], x[277], x[276], x[275], x[274], x[281], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[33], x[292], x[291], x[290], x[289], x[278], x[277], x[276], x[275], x[274], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[317], x[302], x[285], x[316], x[315], x[300], x[282], x[314], x[313], x[298], x[279], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[33], x[264], x[263], x[262], x[273], x[272], x[271], x[305], x[297], x[296], x[295], x[294], x[293], x[289], x[278], x[277], x[276], x[275], x[274]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[317], x[305], x[33], x[264], x[263], x[262], x[273], x[272], x[271], x[302], x[297], x[296], x[295], x[294], x[293], x[285], x[278], x[277], x[276], x[275], x[274]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[316], x[315], x[310], x[309], x[308], x[307], x[306], x[33], x[264], x[263], x[262], x[273], x[272], x[271], x[300], x[297], x[296], x[295], x[294], x[293], x[282], x[278], x[277], x[276], x[275], x[274]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[314], x[313], x[310], x[309], x[308], x[307], x[306], x[33], x[264], x[263], x[262], x[273], x[272], x[271], x[298], x[297], x[296], x[295], x[294], x[293], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[33], x[264], x[263], x[262], x[273], x[272], x[271], x[305], x[297], x[296], x[295], x[294], x[293], x[289], x[278], x[277], x[276], x[275], x[274]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[330], x[315], x[302], x[329], x[328], x[313], x[300], x[327], x[326], x[311], x[298], x[325], x[324], x[323], x[322], x[321], x[320], x[48], x[47], x[46], x[319], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[318], x[310], x[309], x[308], x[307], x[306], x[305], x[297], x[296], x[295], x[294], x[293]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[330], x[318], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[315], x[310], x[309], x[308], x[307], x[306], x[302], x[297], x[296], x[295], x[294], x[293]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[329], x[328], x[324], x[323], x[322], x[321], x[320], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[313], x[310], x[309], x[308], x[307], x[306], x[300], x[297], x[296], x[295], x[294], x[293]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[327], x[326], x[324], x[323], x[322], x[321], x[320], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[311], x[310], x[309], x[308], x[307], x[306], x[298], x[297], x[296], x[295], x[294], x[293]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[325], x[324], x[323], x[322], x[321], x[320], x[48], x[47], x[46], x[319], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[318], x[310], x[309], x[308], x[307], x[306], x[305], x[297], x[296], x[295], x[294], x[293]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[36], x[35], x[34], x[343], x[328], x[315], x[342], x[42], x[41], x[40], x[341], x[326], x[313], x[340], x[39], x[38], x[37], x[339], x[325], x[311], x[338], x[337], x[336], x[335], x[334], x[333], x[45], x[44], x[43], x[332], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[331], x[324], x[323], x[322], x[321], x[320], x[318], x[310], x[309], x[308], x[307], x[306]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[331], x[36], x[35], x[34], x[343], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[328], x[324], x[323], x[322], x[321], x[320], x[315], x[310], x[309], x[308], x[307], x[306]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[342], x[337], x[336], x[335], x[334], x[333], x[42], x[41], x[40], x[341], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[326], x[324], x[323], x[322], x[321], x[320], x[313], x[310], x[309], x[308], x[307], x[306]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[340], x[337], x[336], x[335], x[334], x[333], x[39], x[38], x[37], x[339], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[325], x[324], x[323], x[322], x[321], x[320], x[311], x[310], x[309], x[308], x[307], x[306]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[338], x[337], x[336], x[335], x[334], x[333], x[45], x[44], x[43], x[332], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[331], x[324], x[323], x[322], x[321], x[320], x[318], x[310], x[309], x[308], x[307], x[306]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[356], x[342], x[328], x[355], x[354], x[340], x[326], x[353], x[352], x[338], x[325], x[351], x[350], x[349], x[348], x[347], x[346], x[345], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[344], x[337], x[336], x[335], x[334], x[333], x[331], x[324], x[323], x[322], x[321], x[320]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[356], x[344], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[342], x[337], x[336], x[335], x[334], x[333], x[328], x[324], x[323], x[322], x[321], x[320]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[355], x[354], x[349], x[348], x[347], x[346], x[345], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[340], x[337], x[336], x[335], x[334], x[333], x[326], x[324], x[323], x[322], x[321], x[320]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[353], x[352], x[349], x[348], x[347], x[346], x[345], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[338], x[337], x[336], x[335], x[334], x[333], x[325], x[324], x[323], x[322], x[321], x[320]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[351], x[350], x[349], x[348], x[347], x[346], x[345], x[33], x[264], x[263], x[262], x[51], x[50], x[49], x[344], x[337], x[336], x[335], x[334], x[333], x[331], x[324], x[323], x[322], x[321], x[320]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[369], x[354], x[342], x[368], x[367], x[352], x[340], x[366], x[365], x[350], x[338], x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[357], x[349], x[348], x[347], x[346], x[345], x[344], x[337], x[336], x[335], x[334], x[333]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[369], x[357], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[354], x[349], x[348], x[347], x[346], x[345], x[342], x[337], x[336], x[335], x[334], x[333]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[368], x[367], x[362], x[361], x[360], x[359], x[358], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[352], x[349], x[348], x[347], x[346], x[345], x[340], x[337], x[336], x[335], x[334], x[333]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[366], x[365], x[362], x[361], x[360], x[359], x[358], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[350], x[349], x[348], x[347], x[346], x[345], x[338], x[337], x[336], x[335], x[334], x[333]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[364], x[363], x[362], x[361], x[360], x[359], x[358], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[357], x[349], x[348], x[347], x[346], x[345], x[344], x[337], x[336], x[335], x[334], x[333]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[382], x[367], x[354], x[381], x[380], x[365], x[352], x[379], x[378], x[363], x[350], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[370], x[362], x[361], x[360], x[359], x[358], x[357], x[349], x[348], x[347], x[346], x[345]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[382], x[370], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[367], x[362], x[361], x[360], x[359], x[358], x[354], x[349], x[348], x[347], x[346], x[345]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[381], x[380], x[375], x[374], x[373], x[372], x[371], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[365], x[362], x[361], x[360], x[359], x[358], x[352], x[349], x[348], x[347], x[346], x[345]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[379], x[378], x[375], x[374], x[373], x[372], x[371], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[363], x[362], x[361], x[360], x[359], x[358], x[350], x[349], x[348], x[347], x[346], x[345]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[370], x[362], x[361], x[360], x[359], x[358], x[357], x[349], x[348], x[347], x[346], x[345]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[395], x[380], x[367], x[394], x[393], x[378], x[365], x[392], x[391], x[376], x[363], x[390], x[389], x[388], x[387], x[386], x[385], x[384], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[383], x[375], x[374], x[373], x[372], x[371], x[370], x[362], x[361], x[360], x[359], x[358]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[395], x[383], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[380], x[375], x[374], x[373], x[372], x[371], x[367], x[362], x[361], x[360], x[359], x[358]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[394], x[393], x[388], x[387], x[386], x[385], x[384], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[378], x[375], x[374], x[373], x[372], x[371], x[365], x[362], x[361], x[360], x[359], x[358]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[392], x[391], x[388], x[387], x[386], x[385], x[384], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[376], x[375], x[374], x[373], x[372], x[371], x[363], x[362], x[361], x[360], x[359], x[358]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[390], x[389], x[388], x[387], x[386], x[385], x[384], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[383], x[375], x[374], x[373], x[372], x[371], x[370], x[362], x[361], x[360], x[359], x[358]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[408], x[393], x[380], x[407], x[406], x[391], x[378], x[405], x[404], x[389], x[376], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[396], x[388], x[387], x[386], x[385], x[384], x[383], x[375], x[374], x[373], x[372], x[371]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[408], x[396], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[393], x[388], x[387], x[386], x[385], x[384], x[380], x[375], x[374], x[373], x[372], x[371]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[407], x[406], x[401], x[400], x[399], x[398], x[397], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[391], x[388], x[387], x[386], x[385], x[384], x[378], x[375], x[374], x[373], x[372], x[371]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[405], x[404], x[401], x[400], x[399], x[398], x[397], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[389], x[388], x[387], x[386], x[385], x[384], x[376], x[375], x[374], x[373], x[372], x[371]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[396], x[388], x[387], x[386], x[385], x[384], x[383], x[375], x[374], x[373], x[372], x[371]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[415], x[249], x[184], x[183], x[182], x[181], x[180], x[170], x[178], x[414], x[232], x[234], x[413], x[412], x[258], x[411], x[410], x[161], x[160], x[159], x[158], x[157], x[33], x[256], x[255], x[254], x[409], x[169], x[168], x[167], x[166], x[165], x[253], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[415], x[249], x[184], x[183], x[182], x[181], x[180], x[33], x[256], x[255], x[254], x[170], x[169], x[168], x[167], x[166], x[165], x[178], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[33], x[414], x[258], x[256], x[255], x[254], x[232], x[169], x[168], x[167], x[166], x[165], x[234], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[33], x[413], x[256], x[255], x[254], x[412], x[169], x[168], x[167], x[166], x[165], x[258], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[411], x[410], x[161], x[160], x[159], x[158], x[157], x[33], x[256], x[255], x[254], x[409], x[169], x[168], x[167], x[166], x[165], x[253], x[177], x[176], x[175], x[174], x[173], x[57], x[56], x[55]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[423], x[422], x[209], x[208], x[207], x[206], x[205], x[162], x[170], x[421], x[420], x[202], x[201], x[200], x[199], x[198], x[229], x[232], x[419], x[418], x[194], x[193], x[192], x[191], x[190], x[410], x[412], x[33], x[417], x[111], x[81], x[80], x[79], x[78], x[77], x[256], x[255], x[254], x[416], x[161], x[160], x[159], x[158], x[157], x[409], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[423], x[422], x[209], x[208], x[207], x[206], x[205], x[33], x[256], x[255], x[254], x[162], x[161], x[160], x[159], x[158], x[157], x[170], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[421], x[420], x[202], x[201], x[200], x[199], x[198], x[33], x[256], x[255], x[254], x[229], x[161], x[160], x[159], x[158], x[157], x[232], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[33], x[419], x[418], x[194], x[193], x[192], x[191], x[190], x[256], x[255], x[254], x[410], x[161], x[160], x[159], x[158], x[157], x[412], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[33], x[417], x[111], x[81], x[80], x[79], x[78], x[77], x[256], x[255], x[254], x[416], x[161], x[160], x[159], x[158], x[157], x[409], x[169], x[168], x[167], x[166], x[165], x[57], x[56], x[55]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[428], x[112], x[68], x[67], x[66], x[65], x[64], x[210], x[162], x[427], x[122], x[97], x[96], x[95], x[94], x[93], x[245], x[229], x[426], x[153], x[107], x[106], x[105], x[104], x[103], x[422], x[410], x[425], x[187], x[117], x[116], x[115], x[114], x[113], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[424], x[209], x[208], x[207], x[206], x[205], x[416], x[161], x[160], x[159], x[158], x[157]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[33], x[428], x[112], x[68], x[67], x[66], x[65], x[64], x[57], x[56], x[55], x[256], x[255], x[254], x[210], x[209], x[208], x[207], x[206], x[205], x[162], x[161], x[160], x[159], x[158], x[157]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[33], x[427], x[122], x[97], x[96], x[95], x[94], x[93], x[57], x[56], x[55], x[256], x[255], x[254], x[245], x[209], x[208], x[207], x[206], x[205], x[229], x[161], x[160], x[159], x[158], x[157]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[33], x[426], x[153], x[107], x[106], x[105], x[104], x[103], x[57], x[56], x[55], x[256], x[255], x[254], x[422], x[209], x[208], x[207], x[206], x[205], x[410], x[161], x[160], x[159], x[158], x[157]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[425], x[187], x[117], x[116], x[115], x[114], x[113], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[424], x[209], x[208], x[207], x[206], x[205], x[416], x[161], x[160], x[159], x[158], x[157]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[433], x[212], x[150], x[149], x[148], x[147], x[146], x[203], x[210], x[432], x[219], x[143], x[142], x[141], x[140], x[139], x[243], x[245], x[431], x[228], x[135], x[134], x[133], x[132], x[131], x[420], x[422], x[430], x[238], x[127], x[126], x[125], x[124], x[123], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[429], x[202], x[201], x[200], x[199], x[198], x[424], x[209], x[208], x[207], x[206], x[205]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[433], x[212], x[150], x[149], x[148], x[147], x[146], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[203], x[202], x[201], x[200], x[199], x[198], x[210], x[209], x[208], x[207], x[206], x[205]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[432], x[219], x[143], x[142], x[141], x[140], x[139], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[243], x[202], x[201], x[200], x[199], x[198], x[245], x[209], x[208], x[207], x[206], x[205]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[431], x[228], x[135], x[134], x[133], x[132], x[131], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[420], x[202], x[201], x[200], x[199], x[198], x[422], x[209], x[208], x[207], x[206], x[205]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[430], x[238], x[127], x[126], x[125], x[124], x[123], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[429], x[202], x[201], x[200], x[199], x[198], x[424], x[209], x[208], x[207], x[206], x[205]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[438], x[247], x[184], x[183], x[182], x[181], x[180], x[195], x[203], x[437], x[253], x[177], x[176], x[175], x[174], x[173], x[241], x[243], x[436], x[409], x[169], x[168], x[167], x[166], x[165], x[418], x[420], x[435], x[416], x[161], x[160], x[159], x[158], x[157], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[434], x[194], x[193], x[192], x[191], x[190], x[429], x[202], x[201], x[200], x[199], x[198]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[438], x[247], x[184], x[183], x[182], x[181], x[180], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[195], x[194], x[193], x[192], x[191], x[190], x[203], x[202], x[201], x[200], x[199], x[198]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[437], x[253], x[177], x[176], x[175], x[174], x[173], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[241], x[194], x[193], x[192], x[191], x[190], x[243], x[202], x[201], x[200], x[199], x[198]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[436], x[409], x[169], x[168], x[167], x[166], x[165], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[418], x[194], x[193], x[192], x[191], x[190], x[420], x[202], x[201], x[200], x[199], x[198]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[435], x[416], x[161], x[160], x[159], x[158], x[157], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[434], x[194], x[193], x[192], x[191], x[190], x[429], x[202], x[201], x[200], x[199], x[198]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[442], x[424], x[209], x[208], x[207], x[206], x[205], x[82], x[195], x[441], x[429], x[202], x[201], x[200], x[199], x[198], x[101], x[241], x[440], x[111], x[418], x[33], x[439], x[57], x[56], x[55], x[256], x[255], x[254], x[121], x[81], x[80], x[79], x[78], x[77], x[434], x[194], x[193], x[192], x[191], x[190]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[33], x[442], x[424], x[209], x[208], x[207], x[206], x[205], x[57], x[56], x[55], x[256], x[255], x[254], x[82], x[81], x[80], x[79], x[78], x[77], x[195], x[194], x[193], x[192], x[191], x[190]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[33], x[441], x[429], x[202], x[201], x[200], x[199], x[198], x[57], x[56], x[55], x[256], x[255], x[254], x[101], x[81], x[80], x[79], x[78], x[77], x[241], x[194], x[193], x[192], x[191], x[190]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[440], x[434], x[33], x[57], x[56], x[55], x[256], x[255], x[254], x[111], x[81], x[80], x[79], x[78], x[77], x[418], x[194], x[193], x[192], x[191], x[190]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[33], x[439], x[57], x[56], x[55], x[256], x[255], x[254], x[121], x[81], x[80], x[79], x[78], x[77], x[434], x[194], x[193], x[192], x[191], x[190]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[455], x[406], x[393], x[454], x[453], x[404], x[391], x[452], x[451], x[402], x[389], x[450], x[449], x[448], x[447], x[446], x[445], x[444], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[443], x[401], x[400], x[399], x[398], x[397], x[396], x[388], x[387], x[386], x[385], x[384]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[455], x[443], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[406], x[401], x[400], x[399], x[398], x[397], x[393], x[388], x[387], x[386], x[385], x[384]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[454], x[453], x[448], x[447], x[446], x[445], x[444], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[404], x[401], x[400], x[399], x[398], x[397], x[391], x[388], x[387], x[386], x[385], x[384]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[452], x[451], x[448], x[447], x[446], x[445], x[444], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[402], x[401], x[400], x[399], x[398], x[397], x[389], x[388], x[387], x[386], x[385], x[384]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[450], x[449], x[448], x[447], x[446], x[445], x[444], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[443], x[401], x[400], x[399], x[398], x[397], x[396], x[388], x[387], x[386], x[385], x[384]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[468], x[453], x[406], x[467], x[466], x[451], x[404], x[465], x[464], x[449], x[402], x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[456], x[448], x[447], x[446], x[445], x[444], x[443], x[401], x[400], x[399], x[398], x[397]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[468], x[456], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[453], x[448], x[447], x[446], x[445], x[444], x[406], x[401], x[400], x[399], x[398], x[397]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[467], x[466], x[461], x[460], x[459], x[458], x[457], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[451], x[448], x[447], x[446], x[445], x[444], x[404], x[401], x[400], x[399], x[398], x[397]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[465], x[464], x[461], x[460], x[459], x[458], x[457], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[449], x[448], x[447], x[446], x[445], x[444], x[402], x[401], x[400], x[399], x[398], x[397]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[463], x[462], x[461], x[460], x[459], x[458], x[457], x[33], x[264], x[263], x[262], x[292], x[291], x[290], x[456], x[448], x[447], x[446], x[445], x[444], x[443], x[401], x[400], x[399], x[398], x[397]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[484], x[466], x[453], x[483], x[482], x[464], x[451], x[481], x[480], x[462], x[449], x[479], x[478], x[477], x[476], x[475], x[474], x[473], x[33], x[292], x[291], x[290], x[472], x[461], x[460], x[459], x[458], x[457], x[456], x[448], x[447], x[446], x[445], x[444], x[471], x[470], x[469]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[484], x[472], x[33], x[292], x[291], x[290], x[466], x[461], x[460], x[459], x[458], x[457], x[453], x[448], x[447], x[446], x[445], x[444], x[471], x[470], x[469]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[483], x[482], x[477], x[476], x[475], x[474], x[473], x[33], x[292], x[291], x[290], x[464], x[461], x[460], x[459], x[458], x[457], x[451], x[448], x[447], x[446], x[445], x[444], x[471], x[470], x[469]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[481], x[480], x[477], x[476], x[475], x[474], x[473], x[33], x[292], x[291], x[290], x[462], x[461], x[460], x[459], x[458], x[457], x[449], x[448], x[447], x[446], x[445], x[444], x[471], x[470], x[469]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[479], x[478], x[477], x[476], x[475], x[474], x[473], x[33], x[292], x[291], x[290], x[472], x[461], x[460], x[459], x[458], x[457], x[456], x[448], x[447], x[446], x[445], x[444], x[471], x[470], x[469]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[497], x[482], x[466], x[496], x[495], x[480], x[464], x[494], x[493], x[478], x[462], x[492], x[491], x[490], x[489], x[488], x[487], x[486], x[33], x[273], x[272], x[271], x[485], x[477], x[476], x[475], x[474], x[473], x[472], x[461], x[460], x[459], x[458], x[457], x[471], x[470], x[469]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[497], x[485], x[33], x[273], x[272], x[271], x[482], x[477], x[476], x[475], x[474], x[473], x[466], x[461], x[460], x[459], x[458], x[457], x[471], x[470], x[469]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[496], x[495], x[490], x[489], x[488], x[487], x[486], x[33], x[273], x[272], x[271], x[480], x[477], x[476], x[475], x[474], x[473], x[464], x[461], x[460], x[459], x[458], x[457], x[471], x[470], x[469]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[494], x[493], x[490], x[489], x[488], x[487], x[486], x[33], x[273], x[272], x[271], x[478], x[477], x[476], x[475], x[474], x[473], x[462], x[461], x[460], x[459], x[458], x[457], x[471], x[470], x[469]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[492], x[491], x[490], x[489], x[488], x[487], x[486], x[33], x[273], x[272], x[271], x[485], x[477], x[476], x[475], x[474], x[473], x[472], x[461], x[460], x[459], x[458], x[457], x[471], x[470], x[469]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[510], x[495], x[482], x[509], x[508], x[493], x[480], x[507], x[506], x[491], x[478], x[505], x[504], x[503], x[502], x[501], x[500], x[499], x[33], x[273], x[272], x[271], x[498], x[490], x[489], x[488], x[487], x[486], x[485], x[477], x[476], x[475], x[474], x[473], x[471], x[470], x[469]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[510], x[498], x[33], x[273], x[272], x[271], x[495], x[490], x[489], x[488], x[487], x[486], x[482], x[477], x[476], x[475], x[474], x[473], x[471], x[470], x[469]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[509], x[508], x[503], x[502], x[501], x[500], x[499], x[33], x[273], x[272], x[271], x[493], x[490], x[489], x[488], x[487], x[486], x[480], x[477], x[476], x[475], x[474], x[473], x[471], x[470], x[469]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[507], x[506], x[503], x[502], x[501], x[500], x[499], x[33], x[273], x[272], x[271], x[491], x[490], x[489], x[488], x[487], x[486], x[478], x[477], x[476], x[475], x[474], x[473], x[471], x[470], x[469]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[505], x[504], x[503], x[502], x[501], x[500], x[499], x[33], x[273], x[272], x[271], x[498], x[490], x[489], x[488], x[487], x[486], x[485], x[477], x[476], x[475], x[474], x[473], x[471], x[470], x[469]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[523], x[508], x[495], x[522], x[521], x[506], x[493], x[520], x[519], x[504], x[491], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[511], x[503], x[502], x[501], x[500], x[499], x[498], x[490], x[489], x[488], x[487], x[486]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[523], x[511], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[508], x[503], x[502], x[501], x[500], x[499], x[495], x[490], x[489], x[488], x[487], x[486]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[522], x[521], x[516], x[515], x[514], x[513], x[512], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[506], x[503], x[502], x[501], x[500], x[499], x[493], x[490], x[489], x[488], x[487], x[486]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[520], x[519], x[516], x[515], x[514], x[513], x[512], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[504], x[503], x[502], x[501], x[500], x[499], x[491], x[490], x[489], x[488], x[487], x[486]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[511], x[503], x[502], x[501], x[500], x[499], x[498], x[490], x[489], x[488], x[487], x[486]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[536], x[521], x[508], x[535], x[534], x[519], x[506], x[533], x[532], x[517], x[504], x[531], x[530], x[529], x[528], x[527], x[526], x[525], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[524], x[516], x[515], x[514], x[513], x[512], x[511], x[503], x[502], x[501], x[500], x[499]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[536], x[524], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[521], x[516], x[515], x[514], x[513], x[512], x[508], x[503], x[502], x[501], x[500], x[499]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[535], x[534], x[529], x[528], x[527], x[526], x[525], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[519], x[516], x[515], x[514], x[513], x[512], x[506], x[503], x[502], x[501], x[500], x[499]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[533], x[532], x[529], x[528], x[527], x[526], x[525], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[517], x[516], x[515], x[514], x[513], x[512], x[504], x[503], x[502], x[501], x[500], x[499]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[531], x[530], x[529], x[528], x[527], x[526], x[525], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[524], x[516], x[515], x[514], x[513], x[512], x[511], x[503], x[502], x[501], x[500], x[499]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[549], x[534], x[521], x[548], x[547], x[532], x[519], x[546], x[545], x[530], x[517], x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[537], x[529], x[528], x[527], x[526], x[525], x[524], x[516], x[515], x[514], x[513], x[512]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[549], x[537], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[534], x[529], x[528], x[527], x[526], x[525], x[521], x[516], x[515], x[514], x[513], x[512]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[548], x[547], x[542], x[541], x[540], x[539], x[538], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[532], x[529], x[528], x[527], x[526], x[525], x[519], x[516], x[515], x[514], x[513], x[512]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[546], x[545], x[542], x[541], x[540], x[539], x[538], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[530], x[529], x[528], x[527], x[526], x[525], x[517], x[516], x[515], x[514], x[513], x[512]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[537], x[529], x[528], x[527], x[526], x[525], x[524], x[516], x[515], x[514], x[513], x[512]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[554], x[547], x[534], x[553], x[76], x[545], x[532], x[552], x[100], x[543], x[530], x[551], x[110], x[75], x[74], x[73], x[72], x[71], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[550], x[542], x[541], x[540], x[539], x[538], x[537], x[529], x[528], x[527], x[526], x[525]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[554], x[550], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[547], x[542], x[541], x[540], x[539], x[538], x[534], x[529], x[528], x[527], x[526], x[525]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[553], x[76], x[75], x[74], x[73], x[72], x[71], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[545], x[542], x[541], x[540], x[539], x[538], x[532], x[529], x[528], x[527], x[526], x[525]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[552], x[100], x[75], x[74], x[73], x[72], x[71], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[543], x[542], x[541], x[540], x[539], x[538], x[530], x[529], x[528], x[527], x[526], x[525]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[551], x[110], x[75], x[74], x[73], x[72], x[71], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[550], x[542], x[541], x[540], x[539], x[538], x[537], x[529], x[528], x[527], x[526], x[525]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[558], x[76], x[547], x[557], x[100], x[545], x[556], x[110], x[543], x[91], x[90], x[88], x[89], x[87], x[86], x[85], x[84], x[83], x[555], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[120], x[75], x[74], x[73], x[72], x[71], x[550], x[542], x[541], x[540], x[539], x[538]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[558], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[76], x[75], x[74], x[73], x[72], x[71], x[547], x[542], x[541], x[540], x[539], x[538]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[90], x[91], x[88], x[89], x[87], x[86], x[85], x[84], x[83], x[557], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[100], x[75], x[74], x[73], x[72], x[71], x[545], x[542], x[541], x[540], x[539], x[538]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[90], x[89], x[88], x[91], x[87], x[86], x[85], x[84], x[83], x[556], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[110], x[75], x[74], x[73], x[72], x[71], x[543], x[542], x[541], x[540], x[539], x[538]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[91], x[90], x[88], x[89], x[87], x[86], x[85], x[84], x[83], x[555], x[33], x[471], x[470], x[469], x[273], x[272], x[271], x[120], x[75], x[74], x[73], x[72], x[71], x[550], x[542], x[541], x[540], x[539], x[538]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[121], x[281], x[111], x[110], x[284], x[101], x[100], x[287], x[269], x[268], x[267], x[266], x[265], x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[120], x[75], x[74], x[73], x[72], x[71]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[121], x[81], x[80], x[79], x[78], x[77], x[120], x[75], x[74], x[73], x[72], x[71], x[281], x[269], x[268], x[267], x[266], x[265]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[111], x[81], x[80], x[79], x[78], x[77], x[110], x[75], x[74], x[73], x[72], x[71], x[284], x[269], x[268], x[267], x[266], x[265]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[101], x[81], x[80], x[79], x[78], x[77], x[100], x[75], x[74], x[73], x[72], x[71], x[287], x[269], x[268], x[267], x[266], x[265]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[20], x[19], x[18], x[11], x[10], x[9], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[120], x[75], x[74], x[73], x[72], x[71]}), .y(y[319]));
endmodule

