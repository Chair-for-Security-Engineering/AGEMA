/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [33:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire T1 ;
    wire T2 ;
    wire T3 ;
    wire T4 ;
    wire T5 ;
    wire T6 ;
    wire T7 ;
    wire T8 ;
    wire T9 ;
    wire T10 ;
    wire T11 ;
    wire T12 ;
    wire T13 ;
    wire T14 ;
    wire T15 ;
    wire T16 ;
    wire T17 ;
    wire T18 ;
    wire T19 ;
    wire T20 ;
    wire T21 ;
    wire T22 ;
    wire T23 ;
    wire T24 ;
    wire T25 ;
    wire T26 ;
    wire T27 ;
    wire M1 ;
    wire M2 ;
    wire M3 ;
    wire M4 ;
    wire M5 ;
    wire M6 ;
    wire M7 ;
    wire M8 ;
    wire M9 ;
    wire M10 ;
    wire M11 ;
    wire M12 ;
    wire M13 ;
    wire M14 ;
    wire M15 ;
    wire M16 ;
    wire M17 ;
    wire M18 ;
    wire M19 ;
    wire M20 ;
    wire M21 ;
    wire M22 ;
    wire M23 ;
    wire M24 ;
    wire M25 ;
    wire M26 ;
    wire M27 ;
    wire M28 ;
    wire M29 ;
    wire M30 ;
    wire M31 ;
    wire M32 ;
    wire M33 ;
    wire M34 ;
    wire M35 ;
    wire M36 ;
    wire M37 ;
    wire M38 ;
    wire M39 ;
    wire M40 ;
    wire M41 ;
    wire M42 ;
    wire M43 ;
    wire M44 ;
    wire M45 ;
    wire M46 ;
    wire M47 ;
    wire M48 ;
    wire M49 ;
    wire M50 ;
    wire M51 ;
    wire M52 ;
    wire M53 ;
    wire M54 ;
    wire M55 ;
    wire M56 ;
    wire M57 ;
    wire M58 ;
    wire M59 ;
    wire M60 ;
    wire M61 ;
    wire M62 ;
    wire M63 ;
    wire L0 ;
    wire L1 ;
    wire L2 ;
    wire L3 ;
    wire L4 ;
    wire L5 ;
    wire L6 ;
    wire L7 ;
    wire L8 ;
    wire L9 ;
    wire L10 ;
    wire L11 ;
    wire L12 ;
    wire L13 ;
    wire L14 ;
    wire L15 ;
    wire L16 ;
    wire L17 ;
    wire L18 ;
    wire L19 ;
    wire L20 ;
    wire L21 ;
    wire L22 ;
    wire L23 ;
    wire L24 ;
    wire L25 ;
    wire L26 ;
    wire L27 ;
    wire L28 ;
    wire L29 ;
    wire [7:0] O ;
    wire new_AGEMA_signal_153 ;
    wire new_AGEMA_signal_155 ;
    wire new_AGEMA_signal_157 ;
    wire new_AGEMA_signal_158 ;
    wire new_AGEMA_signal_160 ;
    wire new_AGEMA_signal_163 ;
    wire new_AGEMA_signal_164 ;
    wire new_AGEMA_signal_165 ;
    wire new_AGEMA_signal_167 ;
    wire new_AGEMA_signal_168 ;
    wire new_AGEMA_signal_169 ;
    wire new_AGEMA_signal_170 ;
    wire new_AGEMA_signal_171 ;
    wire new_AGEMA_signal_172 ;
    wire new_AGEMA_signal_173 ;
    wire new_AGEMA_signal_174 ;
    wire new_AGEMA_signal_175 ;
    wire new_AGEMA_signal_176 ;
    wire new_AGEMA_signal_177 ;
    wire new_AGEMA_signal_178 ;
    wire new_AGEMA_signal_179 ;
    wire new_AGEMA_signal_180 ;
    wire new_AGEMA_signal_181 ;
    wire new_AGEMA_signal_182 ;
    wire new_AGEMA_signal_183 ;
    wire new_AGEMA_signal_184 ;
    wire new_AGEMA_signal_185 ;
    wire new_AGEMA_signal_186 ;
    wire new_AGEMA_signal_187 ;
    wire new_AGEMA_signal_188 ;
    wire new_AGEMA_signal_189 ;
    wire new_AGEMA_signal_190 ;
    wire new_AGEMA_signal_191 ;
    wire new_AGEMA_signal_192 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T1_U1 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_153, T1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T2_U1 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_155, T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T3_U1 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_157, T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T4_U1 ( .a ({X_s1[4], X_s0[4]}), .b ({X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_158, T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T5_U1 ( .a ({X_s1[3], X_s0[3]}), .b ({X_s1[1], X_s0[1]}), .c ({new_AGEMA_signal_160, T5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T6_U1 ( .a ({new_AGEMA_signal_153, T1}), .b ({new_AGEMA_signal_160, T5}), .c ({new_AGEMA_signal_169, T6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T7_U1 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[5], X_s0[5]}), .c ({new_AGEMA_signal_163, T7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T8_U1 ( .a ({X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_169, T6}), .c ({new_AGEMA_signal_177, T8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T9_U1 ( .a ({X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_163, T7}), .c ({new_AGEMA_signal_170, T9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T10_U1 ( .a ({new_AGEMA_signal_169, T6}), .b ({new_AGEMA_signal_163, T7}), .c ({new_AGEMA_signal_178, T10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T11_U1 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_164, T11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T12_U1 ( .a ({X_s1[5], X_s0[5]}), .b ({X_s1[2], X_s0[2]}), .c ({new_AGEMA_signal_165, T12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T13_U1 ( .a ({new_AGEMA_signal_157, T3}), .b ({new_AGEMA_signal_158, T4}), .c ({new_AGEMA_signal_171, T13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T14_U1 ( .a ({new_AGEMA_signal_169, T6}), .b ({new_AGEMA_signal_164, T11}), .c ({new_AGEMA_signal_179, T14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T15_U1 ( .a ({new_AGEMA_signal_160, T5}), .b ({new_AGEMA_signal_164, T11}), .c ({new_AGEMA_signal_172, T15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T16_U1 ( .a ({new_AGEMA_signal_160, T5}), .b ({new_AGEMA_signal_165, T12}), .c ({new_AGEMA_signal_173, T16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T17_U1 ( .a ({new_AGEMA_signal_170, T9}), .b ({new_AGEMA_signal_173, T16}), .c ({new_AGEMA_signal_180, T17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T18_U1 ( .a ({X_s1[4], X_s0[4]}), .b ({X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_167, T18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T19_U1 ( .a ({new_AGEMA_signal_163, T7}), .b ({new_AGEMA_signal_167, T18}), .c ({new_AGEMA_signal_174, T19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T20_U1 ( .a ({new_AGEMA_signal_153, T1}), .b ({new_AGEMA_signal_174, T19}), .c ({new_AGEMA_signal_181, T20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T21_U1 ( .a ({X_s1[1], X_s0[1]}), .b ({X_s1[0], X_s0[0]}), .c ({new_AGEMA_signal_168, T21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T22_U1 ( .a ({new_AGEMA_signal_163, T7}), .b ({new_AGEMA_signal_168, T21}), .c ({new_AGEMA_signal_175, T22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T23_U1 ( .a ({new_AGEMA_signal_155, T2}), .b ({new_AGEMA_signal_175, T22}), .c ({new_AGEMA_signal_182, T23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T24_U1 ( .a ({new_AGEMA_signal_155, T2}), .b ({new_AGEMA_signal_178, T10}), .c ({new_AGEMA_signal_190, T24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T25_U1 ( .a ({new_AGEMA_signal_181, T20}), .b ({new_AGEMA_signal_180, T17}), .c ({new_AGEMA_signal_191, T25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T26_U1 ( .a ({new_AGEMA_signal_157, T3}), .b ({new_AGEMA_signal_173, T16}), .c ({new_AGEMA_signal_183, T26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_T27_U1 ( .a ({new_AGEMA_signal_153, T1}), .b ({new_AGEMA_signal_165, T12}), .c ({new_AGEMA_signal_176, T27}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_136 ( .C (clk), .D (T14), .Q (new_AGEMA_signal_329) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C (clk), .D (new_AGEMA_signal_179), .Q (new_AGEMA_signal_331) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C (clk), .D (T26), .Q (new_AGEMA_signal_333) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C (clk), .D (new_AGEMA_signal_183), .Q (new_AGEMA_signal_335) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C (clk), .D (T24), .Q (new_AGEMA_signal_337) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C (clk), .D (new_AGEMA_signal_190), .Q (new_AGEMA_signal_339) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C (clk), .D (T25), .Q (new_AGEMA_signal_341) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C (clk), .D (new_AGEMA_signal_191), .Q (new_AGEMA_signal_343) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C (clk), .D (T6), .Q (new_AGEMA_signal_377) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C (clk), .D (new_AGEMA_signal_169), .Q (new_AGEMA_signal_383) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C (clk), .D (T8), .Q (new_AGEMA_signal_389) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C (clk), .D (new_AGEMA_signal_177), .Q (new_AGEMA_signal_395) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C (clk), .D (X_s0[0]), .Q (new_AGEMA_signal_401) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C (clk), .D (X_s1[0]), .Q (new_AGEMA_signal_407) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C (clk), .D (T16), .Q (new_AGEMA_signal_413) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C (clk), .D (new_AGEMA_signal_173), .Q (new_AGEMA_signal_419) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C (clk), .D (T9), .Q (new_AGEMA_signal_425) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C (clk), .D (new_AGEMA_signal_170), .Q (new_AGEMA_signal_431) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C (clk), .D (T17), .Q (new_AGEMA_signal_437) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C (clk), .D (new_AGEMA_signal_180), .Q (new_AGEMA_signal_443) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C (clk), .D (T15), .Q (new_AGEMA_signal_449) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C (clk), .D (new_AGEMA_signal_172), .Q (new_AGEMA_signal_455) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C (clk), .D (T27), .Q (new_AGEMA_signal_461) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C (clk), .D (new_AGEMA_signal_176), .Q (new_AGEMA_signal_467) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C (clk), .D (T10), .Q (new_AGEMA_signal_473) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C (clk), .D (new_AGEMA_signal_178), .Q (new_AGEMA_signal_479) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C (clk), .D (T13), .Q (new_AGEMA_signal_485) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C (clk), .D (new_AGEMA_signal_171), .Q (new_AGEMA_signal_491) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C (clk), .D (T23), .Q (new_AGEMA_signal_497) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C (clk), .D (new_AGEMA_signal_182), .Q (new_AGEMA_signal_503) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C (clk), .D (T19), .Q (new_AGEMA_signal_509) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C (clk), .D (new_AGEMA_signal_174), .Q (new_AGEMA_signal_515) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C (clk), .D (T3), .Q (new_AGEMA_signal_521) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C (clk), .D (new_AGEMA_signal_157), .Q (new_AGEMA_signal_527) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C (clk), .D (T22), .Q (new_AGEMA_signal_533) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C (clk), .D (new_AGEMA_signal_175), .Q (new_AGEMA_signal_539) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C (clk), .D (T20), .Q (new_AGEMA_signal_545) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C (clk), .D (new_AGEMA_signal_181), .Q (new_AGEMA_signal_551) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C (clk), .D (T1), .Q (new_AGEMA_signal_557) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C (clk), .D (new_AGEMA_signal_153), .Q (new_AGEMA_signal_563) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C (clk), .D (T4), .Q (new_AGEMA_signal_569) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C (clk), .D (new_AGEMA_signal_158), .Q (new_AGEMA_signal_575) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C (clk), .D (T2), .Q (new_AGEMA_signal_581) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C (clk), .D (new_AGEMA_signal_155), .Q (new_AGEMA_signal_587) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M1_U1 ( .a ({new_AGEMA_signal_171, T13}), .b ({new_AGEMA_signal_169, T6}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_184, M1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M2_U1 ( .a ({new_AGEMA_signal_182, T23}), .b ({new_AGEMA_signal_177, T8}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_192, M2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M3_U1 ( .a ({new_AGEMA_signal_332, new_AGEMA_signal_330}), .b ({new_AGEMA_signal_184, M1}), .c ({new_AGEMA_signal_193, M3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M4_U1 ( .a ({new_AGEMA_signal_174, T19}), .b ({X_s1[0], X_s0[0]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_185, M4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M5_U1 ( .a ({new_AGEMA_signal_185, M4}), .b ({new_AGEMA_signal_184, M1}), .c ({new_AGEMA_signal_194, M5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M6_U1 ( .a ({new_AGEMA_signal_157, T3}), .b ({new_AGEMA_signal_173, T16}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_186, M6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M7_U1 ( .a ({new_AGEMA_signal_175, T22}), .b ({new_AGEMA_signal_170, T9}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_187, M7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M8_U1 ( .a ({new_AGEMA_signal_336, new_AGEMA_signal_334}), .b ({new_AGEMA_signal_186, M6}), .c ({new_AGEMA_signal_195, M8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M9_U1 ( .a ({new_AGEMA_signal_181, T20}), .b ({new_AGEMA_signal_180, T17}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_196, M9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M10_U1 ( .a ({new_AGEMA_signal_196, M9}), .b ({new_AGEMA_signal_186, M6}), .c ({new_AGEMA_signal_199, M10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M11_U1 ( .a ({new_AGEMA_signal_153, T1}), .b ({new_AGEMA_signal_172, T15}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_188, M11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M12_U1 ( .a ({new_AGEMA_signal_158, T4}), .b ({new_AGEMA_signal_176, T27}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_189, M12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M13_U1 ( .a ({new_AGEMA_signal_189, M12}), .b ({new_AGEMA_signal_188, M11}), .c ({new_AGEMA_signal_197, M13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M14_U1 ( .a ({new_AGEMA_signal_155, T2}), .b ({new_AGEMA_signal_178, T10}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_198, M14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M15_U1 ( .a ({new_AGEMA_signal_198, M14}), .b ({new_AGEMA_signal_188, M11}), .c ({new_AGEMA_signal_200, M15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M16_U1 ( .a ({new_AGEMA_signal_193, M3}), .b ({new_AGEMA_signal_192, M2}), .c ({new_AGEMA_signal_201, M16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M17_U1 ( .a ({new_AGEMA_signal_194, M5}), .b ({new_AGEMA_signal_340, new_AGEMA_signal_338}), .c ({new_AGEMA_signal_202, M17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M18_U1 ( .a ({new_AGEMA_signal_195, M8}), .b ({new_AGEMA_signal_187, M7}), .c ({new_AGEMA_signal_203, M18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M19_U1 ( .a ({new_AGEMA_signal_199, M10}), .b ({new_AGEMA_signal_200, M15}), .c ({new_AGEMA_signal_204, M19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M20_U1 ( .a ({new_AGEMA_signal_201, M16}), .b ({new_AGEMA_signal_197, M13}), .c ({new_AGEMA_signal_205, M20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M21_U1 ( .a ({new_AGEMA_signal_202, M17}), .b ({new_AGEMA_signal_200, M15}), .c ({new_AGEMA_signal_206, M21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M22_U1 ( .a ({new_AGEMA_signal_203, M18}), .b ({new_AGEMA_signal_197, M13}), .c ({new_AGEMA_signal_207, M22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M23_U1 ( .a ({new_AGEMA_signal_204, M19}), .b ({new_AGEMA_signal_344, new_AGEMA_signal_342}), .c ({new_AGEMA_signal_208, M23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M24_U1 ( .a ({new_AGEMA_signal_207, M22}), .b ({new_AGEMA_signal_208, M23}), .c ({new_AGEMA_signal_212, M24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M27_U1 ( .a ({new_AGEMA_signal_205, M20}), .b ({new_AGEMA_signal_206, M21}), .c ({new_AGEMA_signal_210, M27}) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C (clk), .D (new_AGEMA_signal_329), .Q (new_AGEMA_signal_330) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C (clk), .D (new_AGEMA_signal_331), .Q (new_AGEMA_signal_332) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C (clk), .D (new_AGEMA_signal_333), .Q (new_AGEMA_signal_334) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C (clk), .D (new_AGEMA_signal_335), .Q (new_AGEMA_signal_336) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C (clk), .D (new_AGEMA_signal_337), .Q (new_AGEMA_signal_338) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C (clk), .D (new_AGEMA_signal_339), .Q (new_AGEMA_signal_340) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C (clk), .D (new_AGEMA_signal_341), .Q (new_AGEMA_signal_342) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C (clk), .D (new_AGEMA_signal_343), .Q (new_AGEMA_signal_344) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C (clk), .D (new_AGEMA_signal_377), .Q (new_AGEMA_signal_378) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C (clk), .D (new_AGEMA_signal_383), .Q (new_AGEMA_signal_384) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C (clk), .D (new_AGEMA_signal_389), .Q (new_AGEMA_signal_390) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C (clk), .D (new_AGEMA_signal_395), .Q (new_AGEMA_signal_396) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C (clk), .D (new_AGEMA_signal_401), .Q (new_AGEMA_signal_402) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C (clk), .D (new_AGEMA_signal_407), .Q (new_AGEMA_signal_408) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C (clk), .D (new_AGEMA_signal_413), .Q (new_AGEMA_signal_414) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C (clk), .D (new_AGEMA_signal_419), .Q (new_AGEMA_signal_420) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C (clk), .D (new_AGEMA_signal_425), .Q (new_AGEMA_signal_426) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C (clk), .D (new_AGEMA_signal_431), .Q (new_AGEMA_signal_432) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C (clk), .D (new_AGEMA_signal_437), .Q (new_AGEMA_signal_438) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C (clk), .D (new_AGEMA_signal_443), .Q (new_AGEMA_signal_444) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C (clk), .D (new_AGEMA_signal_449), .Q (new_AGEMA_signal_450) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C (clk), .D (new_AGEMA_signal_455), .Q (new_AGEMA_signal_456) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C (clk), .D (new_AGEMA_signal_461), .Q (new_AGEMA_signal_462) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C (clk), .D (new_AGEMA_signal_467), .Q (new_AGEMA_signal_468) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C (clk), .D (new_AGEMA_signal_473), .Q (new_AGEMA_signal_474) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C (clk), .D (new_AGEMA_signal_479), .Q (new_AGEMA_signal_480) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C (clk), .D (new_AGEMA_signal_485), .Q (new_AGEMA_signal_486) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C (clk), .D (new_AGEMA_signal_491), .Q (new_AGEMA_signal_492) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C (clk), .D (new_AGEMA_signal_497), .Q (new_AGEMA_signal_498) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C (clk), .D (new_AGEMA_signal_503), .Q (new_AGEMA_signal_504) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C (clk), .D (new_AGEMA_signal_509), .Q (new_AGEMA_signal_510) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C (clk), .D (new_AGEMA_signal_515), .Q (new_AGEMA_signal_516) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C (clk), .D (new_AGEMA_signal_521), .Q (new_AGEMA_signal_522) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C (clk), .D (new_AGEMA_signal_527), .Q (new_AGEMA_signal_528) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C (clk), .D (new_AGEMA_signal_533), .Q (new_AGEMA_signal_534) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C (clk), .D (new_AGEMA_signal_539), .Q (new_AGEMA_signal_540) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C (clk), .D (new_AGEMA_signal_545), .Q (new_AGEMA_signal_546) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C (clk), .D (new_AGEMA_signal_551), .Q (new_AGEMA_signal_552) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C (clk), .D (new_AGEMA_signal_557), .Q (new_AGEMA_signal_558) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C (clk), .D (new_AGEMA_signal_563), .Q (new_AGEMA_signal_564) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C (clk), .D (new_AGEMA_signal_569), .Q (new_AGEMA_signal_570) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C (clk), .D (new_AGEMA_signal_575), .Q (new_AGEMA_signal_576) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C (clk), .D (new_AGEMA_signal_581), .Q (new_AGEMA_signal_582) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C (clk), .D (new_AGEMA_signal_587), .Q (new_AGEMA_signal_588) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_152 ( .C (clk), .D (M21), .Q (new_AGEMA_signal_345) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C (clk), .D (new_AGEMA_signal_206), .Q (new_AGEMA_signal_347) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C (clk), .D (M23), .Q (new_AGEMA_signal_349) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C (clk), .D (new_AGEMA_signal_208), .Q (new_AGEMA_signal_351) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C (clk), .D (M27), .Q (new_AGEMA_signal_353) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C (clk), .D (new_AGEMA_signal_210), .Q (new_AGEMA_signal_355) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C (clk), .D (M24), .Q (new_AGEMA_signal_357) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C (clk), .D (new_AGEMA_signal_212), .Q (new_AGEMA_signal_359) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C (clk), .D (new_AGEMA_signal_378), .Q (new_AGEMA_signal_379) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C (clk), .D (new_AGEMA_signal_384), .Q (new_AGEMA_signal_385) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C (clk), .D (new_AGEMA_signal_390), .Q (new_AGEMA_signal_391) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C (clk), .D (new_AGEMA_signal_396), .Q (new_AGEMA_signal_397) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C (clk), .D (new_AGEMA_signal_402), .Q (new_AGEMA_signal_403) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C (clk), .D (new_AGEMA_signal_408), .Q (new_AGEMA_signal_409) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C (clk), .D (new_AGEMA_signal_414), .Q (new_AGEMA_signal_415) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C (clk), .D (new_AGEMA_signal_420), .Q (new_AGEMA_signal_421) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C (clk), .D (new_AGEMA_signal_426), .Q (new_AGEMA_signal_427) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C (clk), .D (new_AGEMA_signal_432), .Q (new_AGEMA_signal_433) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C (clk), .D (new_AGEMA_signal_438), .Q (new_AGEMA_signal_439) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C (clk), .D (new_AGEMA_signal_444), .Q (new_AGEMA_signal_445) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C (clk), .D (new_AGEMA_signal_450), .Q (new_AGEMA_signal_451) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C (clk), .D (new_AGEMA_signal_456), .Q (new_AGEMA_signal_457) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C (clk), .D (new_AGEMA_signal_462), .Q (new_AGEMA_signal_463) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C (clk), .D (new_AGEMA_signal_468), .Q (new_AGEMA_signal_469) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C (clk), .D (new_AGEMA_signal_474), .Q (new_AGEMA_signal_475) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C (clk), .D (new_AGEMA_signal_480), .Q (new_AGEMA_signal_481) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C (clk), .D (new_AGEMA_signal_486), .Q (new_AGEMA_signal_487) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C (clk), .D (new_AGEMA_signal_492), .Q (new_AGEMA_signal_493) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C (clk), .D (new_AGEMA_signal_498), .Q (new_AGEMA_signal_499) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C (clk), .D (new_AGEMA_signal_504), .Q (new_AGEMA_signal_505) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C (clk), .D (new_AGEMA_signal_510), .Q (new_AGEMA_signal_511) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C (clk), .D (new_AGEMA_signal_516), .Q (new_AGEMA_signal_517) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C (clk), .D (new_AGEMA_signal_522), .Q (new_AGEMA_signal_523) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C (clk), .D (new_AGEMA_signal_528), .Q (new_AGEMA_signal_529) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C (clk), .D (new_AGEMA_signal_534), .Q (new_AGEMA_signal_535) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C (clk), .D (new_AGEMA_signal_540), .Q (new_AGEMA_signal_541) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C (clk), .D (new_AGEMA_signal_546), .Q (new_AGEMA_signal_547) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C (clk), .D (new_AGEMA_signal_552), .Q (new_AGEMA_signal_553) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C (clk), .D (new_AGEMA_signal_558), .Q (new_AGEMA_signal_559) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C (clk), .D (new_AGEMA_signal_564), .Q (new_AGEMA_signal_565) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C (clk), .D (new_AGEMA_signal_570), .Q (new_AGEMA_signal_571) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C (clk), .D (new_AGEMA_signal_576), .Q (new_AGEMA_signal_577) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C (clk), .D (new_AGEMA_signal_582), .Q (new_AGEMA_signal_583) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C (clk), .D (new_AGEMA_signal_588), .Q (new_AGEMA_signal_589) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M25_U1 ( .a ({new_AGEMA_signal_207, M22}), .b ({new_AGEMA_signal_205, M20}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_209, M25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M26_U1 ( .a ({new_AGEMA_signal_348, new_AGEMA_signal_346}), .b ({new_AGEMA_signal_209, M25}), .c ({new_AGEMA_signal_213, M26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M28_U1 ( .a ({new_AGEMA_signal_352, new_AGEMA_signal_350}), .b ({new_AGEMA_signal_209, M25}), .c ({new_AGEMA_signal_214, M28}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M31_U1 ( .a ({new_AGEMA_signal_205, M20}), .b ({new_AGEMA_signal_208, M23}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_215, M31}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M33_U1 ( .a ({new_AGEMA_signal_356, new_AGEMA_signal_354}), .b ({new_AGEMA_signal_209, M25}), .c ({new_AGEMA_signal_216, M33}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M34_U1 ( .a ({new_AGEMA_signal_206, M21}), .b ({new_AGEMA_signal_207, M22}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_211, M34}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M36_U1 ( .a ({new_AGEMA_signal_360, new_AGEMA_signal_358}), .b ({new_AGEMA_signal_209, M25}), .c ({new_AGEMA_signal_221, M36}) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C (clk), .D (new_AGEMA_signal_345), .Q (new_AGEMA_signal_346) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C (clk), .D (new_AGEMA_signal_347), .Q (new_AGEMA_signal_348) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C (clk), .D (new_AGEMA_signal_349), .Q (new_AGEMA_signal_350) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C (clk), .D (new_AGEMA_signal_351), .Q (new_AGEMA_signal_352) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C (clk), .D (new_AGEMA_signal_353), .Q (new_AGEMA_signal_354) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C (clk), .D (new_AGEMA_signal_355), .Q (new_AGEMA_signal_356) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C (clk), .D (new_AGEMA_signal_357), .Q (new_AGEMA_signal_358) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C (clk), .D (new_AGEMA_signal_359), .Q (new_AGEMA_signal_360) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C (clk), .D (new_AGEMA_signal_379), .Q (new_AGEMA_signal_380) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C (clk), .D (new_AGEMA_signal_385), .Q (new_AGEMA_signal_386) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C (clk), .D (new_AGEMA_signal_391), .Q (new_AGEMA_signal_392) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C (clk), .D (new_AGEMA_signal_397), .Q (new_AGEMA_signal_398) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C (clk), .D (new_AGEMA_signal_403), .Q (new_AGEMA_signal_404) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C (clk), .D (new_AGEMA_signal_409), .Q (new_AGEMA_signal_410) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C (clk), .D (new_AGEMA_signal_415), .Q (new_AGEMA_signal_416) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C (clk), .D (new_AGEMA_signal_421), .Q (new_AGEMA_signal_422) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C (clk), .D (new_AGEMA_signal_427), .Q (new_AGEMA_signal_428) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C (clk), .D (new_AGEMA_signal_433), .Q (new_AGEMA_signal_434) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C (clk), .D (new_AGEMA_signal_439), .Q (new_AGEMA_signal_440) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C (clk), .D (new_AGEMA_signal_445), .Q (new_AGEMA_signal_446) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C (clk), .D (new_AGEMA_signal_451), .Q (new_AGEMA_signal_452) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C (clk), .D (new_AGEMA_signal_457), .Q (new_AGEMA_signal_458) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C (clk), .D (new_AGEMA_signal_463), .Q (new_AGEMA_signal_464) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C (clk), .D (new_AGEMA_signal_469), .Q (new_AGEMA_signal_470) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C (clk), .D (new_AGEMA_signal_475), .Q (new_AGEMA_signal_476) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C (clk), .D (new_AGEMA_signal_481), .Q (new_AGEMA_signal_482) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C (clk), .D (new_AGEMA_signal_487), .Q (new_AGEMA_signal_488) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C (clk), .D (new_AGEMA_signal_493), .Q (new_AGEMA_signal_494) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C (clk), .D (new_AGEMA_signal_499), .Q (new_AGEMA_signal_500) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C (clk), .D (new_AGEMA_signal_505), .Q (new_AGEMA_signal_506) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C (clk), .D (new_AGEMA_signal_511), .Q (new_AGEMA_signal_512) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C (clk), .D (new_AGEMA_signal_517), .Q (new_AGEMA_signal_518) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C (clk), .D (new_AGEMA_signal_523), .Q (new_AGEMA_signal_524) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C (clk), .D (new_AGEMA_signal_529), .Q (new_AGEMA_signal_530) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C (clk), .D (new_AGEMA_signal_535), .Q (new_AGEMA_signal_536) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C (clk), .D (new_AGEMA_signal_541), .Q (new_AGEMA_signal_542) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C (clk), .D (new_AGEMA_signal_547), .Q (new_AGEMA_signal_548) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C (clk), .D (new_AGEMA_signal_553), .Q (new_AGEMA_signal_554) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C (clk), .D (new_AGEMA_signal_559), .Q (new_AGEMA_signal_560) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C (clk), .D (new_AGEMA_signal_565), .Q (new_AGEMA_signal_566) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C (clk), .D (new_AGEMA_signal_571), .Q (new_AGEMA_signal_572) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C (clk), .D (new_AGEMA_signal_577), .Q (new_AGEMA_signal_578) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C (clk), .D (new_AGEMA_signal_583), .Q (new_AGEMA_signal_584) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C (clk), .D (new_AGEMA_signal_589), .Q (new_AGEMA_signal_590) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_168 ( .C (clk), .D (new_AGEMA_signal_346), .Q (new_AGEMA_signal_361) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C (clk), .D (new_AGEMA_signal_348), .Q (new_AGEMA_signal_363) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C (clk), .D (M33), .Q (new_AGEMA_signal_365) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C (clk), .D (new_AGEMA_signal_216), .Q (new_AGEMA_signal_367) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C (clk), .D (new_AGEMA_signal_350), .Q (new_AGEMA_signal_369) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C (clk), .D (new_AGEMA_signal_352), .Q (new_AGEMA_signal_371) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C (clk), .D (M36), .Q (new_AGEMA_signal_373) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C (clk), .D (new_AGEMA_signal_221), .Q (new_AGEMA_signal_375) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C (clk), .D (new_AGEMA_signal_380), .Q (new_AGEMA_signal_381) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C (clk), .D (new_AGEMA_signal_386), .Q (new_AGEMA_signal_387) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C (clk), .D (new_AGEMA_signal_392), .Q (new_AGEMA_signal_393) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C (clk), .D (new_AGEMA_signal_398), .Q (new_AGEMA_signal_399) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C (clk), .D (new_AGEMA_signal_404), .Q (new_AGEMA_signal_405) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C (clk), .D (new_AGEMA_signal_410), .Q (new_AGEMA_signal_411) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C (clk), .D (new_AGEMA_signal_416), .Q (new_AGEMA_signal_417) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C (clk), .D (new_AGEMA_signal_422), .Q (new_AGEMA_signal_423) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C (clk), .D (new_AGEMA_signal_428), .Q (new_AGEMA_signal_429) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C (clk), .D (new_AGEMA_signal_434), .Q (new_AGEMA_signal_435) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C (clk), .D (new_AGEMA_signal_440), .Q (new_AGEMA_signal_441) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C (clk), .D (new_AGEMA_signal_446), .Q (new_AGEMA_signal_447) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C (clk), .D (new_AGEMA_signal_452), .Q (new_AGEMA_signal_453) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C (clk), .D (new_AGEMA_signal_458), .Q (new_AGEMA_signal_459) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C (clk), .D (new_AGEMA_signal_464), .Q (new_AGEMA_signal_465) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C (clk), .D (new_AGEMA_signal_470), .Q (new_AGEMA_signal_471) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C (clk), .D (new_AGEMA_signal_476), .Q (new_AGEMA_signal_477) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C (clk), .D (new_AGEMA_signal_482), .Q (new_AGEMA_signal_483) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C (clk), .D (new_AGEMA_signal_488), .Q (new_AGEMA_signal_489) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C (clk), .D (new_AGEMA_signal_494), .Q (new_AGEMA_signal_495) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C (clk), .D (new_AGEMA_signal_500), .Q (new_AGEMA_signal_501) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C (clk), .D (new_AGEMA_signal_506), .Q (new_AGEMA_signal_507) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C (clk), .D (new_AGEMA_signal_512), .Q (new_AGEMA_signal_513) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C (clk), .D (new_AGEMA_signal_518), .Q (new_AGEMA_signal_519) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C (clk), .D (new_AGEMA_signal_524), .Q (new_AGEMA_signal_525) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C (clk), .D (new_AGEMA_signal_530), .Q (new_AGEMA_signal_531) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C (clk), .D (new_AGEMA_signal_536), .Q (new_AGEMA_signal_537) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C (clk), .D (new_AGEMA_signal_542), .Q (new_AGEMA_signal_543) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C (clk), .D (new_AGEMA_signal_548), .Q (new_AGEMA_signal_549) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C (clk), .D (new_AGEMA_signal_554), .Q (new_AGEMA_signal_555) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C (clk), .D (new_AGEMA_signal_560), .Q (new_AGEMA_signal_561) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C (clk), .D (new_AGEMA_signal_566), .Q (new_AGEMA_signal_567) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C (clk), .D (new_AGEMA_signal_572), .Q (new_AGEMA_signal_573) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C (clk), .D (new_AGEMA_signal_578), .Q (new_AGEMA_signal_579) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C (clk), .D (new_AGEMA_signal_584), .Q (new_AGEMA_signal_585) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C (clk), .D (new_AGEMA_signal_590), .Q (new_AGEMA_signal_591) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M29_U1 ( .a ({new_AGEMA_signal_214, M28}), .b ({new_AGEMA_signal_356, new_AGEMA_signal_354}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_217, M29}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M30_U1 ( .a ({new_AGEMA_signal_213, M26}), .b ({new_AGEMA_signal_360, new_AGEMA_signal_358}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_218, M30}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M32_U1 ( .a ({new_AGEMA_signal_356, new_AGEMA_signal_354}), .b ({new_AGEMA_signal_215, M31}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_219, M32}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M35_U1 ( .a ({new_AGEMA_signal_360, new_AGEMA_signal_358}), .b ({new_AGEMA_signal_211, M34}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_220, M35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M37_U1 ( .a ({new_AGEMA_signal_364, new_AGEMA_signal_362}), .b ({new_AGEMA_signal_217, M29}), .c ({new_AGEMA_signal_222, M37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M38_U1 ( .a ({new_AGEMA_signal_219, M32}), .b ({new_AGEMA_signal_368, new_AGEMA_signal_366}), .c ({new_AGEMA_signal_223, M38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M39_U1 ( .a ({new_AGEMA_signal_372, new_AGEMA_signal_370}), .b ({new_AGEMA_signal_218, M30}), .c ({new_AGEMA_signal_224, M39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M40_U1 ( .a ({new_AGEMA_signal_220, M35}), .b ({new_AGEMA_signal_376, new_AGEMA_signal_374}), .c ({new_AGEMA_signal_225, M40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M41_U1 ( .a ({new_AGEMA_signal_223, M38}), .b ({new_AGEMA_signal_225, M40}), .c ({new_AGEMA_signal_226, M41}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M42_U1 ( .a ({new_AGEMA_signal_222, M37}), .b ({new_AGEMA_signal_224, M39}), .c ({new_AGEMA_signal_227, M42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M43_U1 ( .a ({new_AGEMA_signal_222, M37}), .b ({new_AGEMA_signal_223, M38}), .c ({new_AGEMA_signal_228, M43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M44_U1 ( .a ({new_AGEMA_signal_224, M39}), .b ({new_AGEMA_signal_225, M40}), .c ({new_AGEMA_signal_229, M44}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_M45_U1 ( .a ({new_AGEMA_signal_227, M42}), .b ({new_AGEMA_signal_226, M41}), .c ({new_AGEMA_signal_238, M45}) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C (clk), .D (new_AGEMA_signal_361), .Q (new_AGEMA_signal_362) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C (clk), .D (new_AGEMA_signal_363), .Q (new_AGEMA_signal_364) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C (clk), .D (new_AGEMA_signal_365), .Q (new_AGEMA_signal_366) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C (clk), .D (new_AGEMA_signal_367), .Q (new_AGEMA_signal_368) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C (clk), .D (new_AGEMA_signal_369), .Q (new_AGEMA_signal_370) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C (clk), .D (new_AGEMA_signal_371), .Q (new_AGEMA_signal_372) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C (clk), .D (new_AGEMA_signal_373), .Q (new_AGEMA_signal_374) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C (clk), .D (new_AGEMA_signal_375), .Q (new_AGEMA_signal_376) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C (clk), .D (new_AGEMA_signal_381), .Q (new_AGEMA_signal_382) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C (clk), .D (new_AGEMA_signal_387), .Q (new_AGEMA_signal_388) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C (clk), .D (new_AGEMA_signal_393), .Q (new_AGEMA_signal_394) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C (clk), .D (new_AGEMA_signal_399), .Q (new_AGEMA_signal_400) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C (clk), .D (new_AGEMA_signal_405), .Q (new_AGEMA_signal_406) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C (clk), .D (new_AGEMA_signal_411), .Q (new_AGEMA_signal_412) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C (clk), .D (new_AGEMA_signal_417), .Q (new_AGEMA_signal_418) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C (clk), .D (new_AGEMA_signal_423), .Q (new_AGEMA_signal_424) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C (clk), .D (new_AGEMA_signal_429), .Q (new_AGEMA_signal_430) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C (clk), .D (new_AGEMA_signal_435), .Q (new_AGEMA_signal_436) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C (clk), .D (new_AGEMA_signal_441), .Q (new_AGEMA_signal_442) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C (clk), .D (new_AGEMA_signal_447), .Q (new_AGEMA_signal_448) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C (clk), .D (new_AGEMA_signal_453), .Q (new_AGEMA_signal_454) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C (clk), .D (new_AGEMA_signal_459), .Q (new_AGEMA_signal_460) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C (clk), .D (new_AGEMA_signal_465), .Q (new_AGEMA_signal_466) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C (clk), .D (new_AGEMA_signal_471), .Q (new_AGEMA_signal_472) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C (clk), .D (new_AGEMA_signal_477), .Q (new_AGEMA_signal_478) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C (clk), .D (new_AGEMA_signal_483), .Q (new_AGEMA_signal_484) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C (clk), .D (new_AGEMA_signal_489), .Q (new_AGEMA_signal_490) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C (clk), .D (new_AGEMA_signal_495), .Q (new_AGEMA_signal_496) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C (clk), .D (new_AGEMA_signal_501), .Q (new_AGEMA_signal_502) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C (clk), .D (new_AGEMA_signal_507), .Q (new_AGEMA_signal_508) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C (clk), .D (new_AGEMA_signal_513), .Q (new_AGEMA_signal_514) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C (clk), .D (new_AGEMA_signal_519), .Q (new_AGEMA_signal_520) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C (clk), .D (new_AGEMA_signal_525), .Q (new_AGEMA_signal_526) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C (clk), .D (new_AGEMA_signal_531), .Q (new_AGEMA_signal_532) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C (clk), .D (new_AGEMA_signal_537), .Q (new_AGEMA_signal_538) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C (clk), .D (new_AGEMA_signal_543), .Q (new_AGEMA_signal_544) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C (clk), .D (new_AGEMA_signal_549), .Q (new_AGEMA_signal_550) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C (clk), .D (new_AGEMA_signal_555), .Q (new_AGEMA_signal_556) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C (clk), .D (new_AGEMA_signal_561), .Q (new_AGEMA_signal_562) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C (clk), .D (new_AGEMA_signal_567), .Q (new_AGEMA_signal_568) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C (clk), .D (new_AGEMA_signal_573), .Q (new_AGEMA_signal_574) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C (clk), .D (new_AGEMA_signal_579), .Q (new_AGEMA_signal_580) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C (clk), .D (new_AGEMA_signal_585), .Q (new_AGEMA_signal_586) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C (clk), .D (new_AGEMA_signal_591), .Q (new_AGEMA_signal_592) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M46_U1 ( .a ({new_AGEMA_signal_229, M44}), .b ({new_AGEMA_signal_388, new_AGEMA_signal_382}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_239, M46}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M47_U1 ( .a ({new_AGEMA_signal_225, M40}), .b ({new_AGEMA_signal_400, new_AGEMA_signal_394}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_230, M47}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M48_U1 ( .a ({new_AGEMA_signal_224, M39}), .b ({new_AGEMA_signal_412, new_AGEMA_signal_406}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_231, M48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M49_U1 ( .a ({new_AGEMA_signal_228, M43}), .b ({new_AGEMA_signal_424, new_AGEMA_signal_418}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_240, M49}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M50_U1 ( .a ({new_AGEMA_signal_223, M38}), .b ({new_AGEMA_signal_436, new_AGEMA_signal_430}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_232, M50}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M51_U1 ( .a ({new_AGEMA_signal_222, M37}), .b ({new_AGEMA_signal_448, new_AGEMA_signal_442}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_233, M51}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M52_U1 ( .a ({new_AGEMA_signal_227, M42}), .b ({new_AGEMA_signal_460, new_AGEMA_signal_454}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_241, M52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M53_U1 ( .a ({new_AGEMA_signal_238, M45}), .b ({new_AGEMA_signal_472, new_AGEMA_signal_466}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_250, M53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M54_U1 ( .a ({new_AGEMA_signal_226, M41}), .b ({new_AGEMA_signal_484, new_AGEMA_signal_478}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_242, M54}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M55_U1 ( .a ({new_AGEMA_signal_229, M44}), .b ({new_AGEMA_signal_496, new_AGEMA_signal_490}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_243, M55}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M56_U1 ( .a ({new_AGEMA_signal_225, M40}), .b ({new_AGEMA_signal_508, new_AGEMA_signal_502}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_234, M56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M57_U1 ( .a ({new_AGEMA_signal_224, M39}), .b ({new_AGEMA_signal_520, new_AGEMA_signal_514}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_235, M57}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M58_U1 ( .a ({new_AGEMA_signal_228, M43}), .b ({new_AGEMA_signal_532, new_AGEMA_signal_526}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_244, M58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M59_U1 ( .a ({new_AGEMA_signal_223, M38}), .b ({new_AGEMA_signal_544, new_AGEMA_signal_538}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_236, M59}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M60_U1 ( .a ({new_AGEMA_signal_222, M37}), .b ({new_AGEMA_signal_556, new_AGEMA_signal_550}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_237, M60}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M61_U1 ( .a ({new_AGEMA_signal_227, M42}), .b ({new_AGEMA_signal_568, new_AGEMA_signal_562}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_245, M61}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M62_U1 ( .a ({new_AGEMA_signal_238, M45}), .b ({new_AGEMA_signal_580, new_AGEMA_signal_574}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_251, M62}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) AND_M63_U1 ( .a ({new_AGEMA_signal_226, M41}), .b ({new_AGEMA_signal_592, new_AGEMA_signal_586}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_246, M63}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L0_U1 ( .a ({new_AGEMA_signal_245, M61}), .b ({new_AGEMA_signal_251, M62}), .c ({new_AGEMA_signal_260, L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L1_U1 ( .a ({new_AGEMA_signal_232, M50}), .b ({new_AGEMA_signal_234, M56}), .c ({new_AGEMA_signal_247, L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L2_U1 ( .a ({new_AGEMA_signal_239, M46}), .b ({new_AGEMA_signal_231, M48}), .c ({new_AGEMA_signal_252, L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L3_U1 ( .a ({new_AGEMA_signal_230, M47}), .b ({new_AGEMA_signal_243, M55}), .c ({new_AGEMA_signal_253, L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L4_U1 ( .a ({new_AGEMA_signal_242, M54}), .b ({new_AGEMA_signal_244, M58}), .c ({new_AGEMA_signal_254, L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L5_U1 ( .a ({new_AGEMA_signal_240, M49}), .b ({new_AGEMA_signal_245, M61}), .c ({new_AGEMA_signal_255, L5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L6_U1 ( .a ({new_AGEMA_signal_251, M62}), .b ({new_AGEMA_signal_255, L5}), .c ({new_AGEMA_signal_261, L6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L7_U1 ( .a ({new_AGEMA_signal_239, M46}), .b ({new_AGEMA_signal_253, L3}), .c ({new_AGEMA_signal_262, L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L8_U1 ( .a ({new_AGEMA_signal_233, M51}), .b ({new_AGEMA_signal_236, M59}), .c ({new_AGEMA_signal_248, L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L9_U1 ( .a ({new_AGEMA_signal_241, M52}), .b ({new_AGEMA_signal_250, M53}), .c ({new_AGEMA_signal_263, L9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L10_U1 ( .a ({new_AGEMA_signal_250, M53}), .b ({new_AGEMA_signal_254, L4}), .c ({new_AGEMA_signal_264, L10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L11_U1 ( .a ({new_AGEMA_signal_237, M60}), .b ({new_AGEMA_signal_252, L2}), .c ({new_AGEMA_signal_265, L11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L12_U1 ( .a ({new_AGEMA_signal_231, M48}), .b ({new_AGEMA_signal_233, M51}), .c ({new_AGEMA_signal_249, L12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L13_U1 ( .a ({new_AGEMA_signal_232, M50}), .b ({new_AGEMA_signal_260, L0}), .c ({new_AGEMA_signal_269, L13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L14_U1 ( .a ({new_AGEMA_signal_241, M52}), .b ({new_AGEMA_signal_245, M61}), .c ({new_AGEMA_signal_256, L14}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L15_U1 ( .a ({new_AGEMA_signal_243, M55}), .b ({new_AGEMA_signal_247, L1}), .c ({new_AGEMA_signal_257, L15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L16_U1 ( .a ({new_AGEMA_signal_234, M56}), .b ({new_AGEMA_signal_260, L0}), .c ({new_AGEMA_signal_270, L16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L17_U1 ( .a ({new_AGEMA_signal_235, M57}), .b ({new_AGEMA_signal_247, L1}), .c ({new_AGEMA_signal_258, L17}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L18_U1 ( .a ({new_AGEMA_signal_244, M58}), .b ({new_AGEMA_signal_248, L8}), .c ({new_AGEMA_signal_259, L18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L19_U1 ( .a ({new_AGEMA_signal_246, M63}), .b ({new_AGEMA_signal_254, L4}), .c ({new_AGEMA_signal_266, L19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L20_U1 ( .a ({new_AGEMA_signal_260, L0}), .b ({new_AGEMA_signal_247, L1}), .c ({new_AGEMA_signal_271, L20}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L21_U1 ( .a ({new_AGEMA_signal_247, L1}), .b ({new_AGEMA_signal_262, L7}), .c ({new_AGEMA_signal_272, L21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L22_U1 ( .a ({new_AGEMA_signal_253, L3}), .b ({new_AGEMA_signal_249, L12}), .c ({new_AGEMA_signal_267, L22}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L23_U1 ( .a ({new_AGEMA_signal_259, L18}), .b ({new_AGEMA_signal_252, L2}), .c ({new_AGEMA_signal_268, L23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L24_U1 ( .a ({new_AGEMA_signal_257, L15}), .b ({new_AGEMA_signal_263, L9}), .c ({new_AGEMA_signal_273, L24}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L25_U1 ( .a ({new_AGEMA_signal_261, L6}), .b ({new_AGEMA_signal_264, L10}), .c ({new_AGEMA_signal_274, L25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L26_U1 ( .a ({new_AGEMA_signal_262, L7}), .b ({new_AGEMA_signal_263, L9}), .c ({new_AGEMA_signal_275, L26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L27_U1 ( .a ({new_AGEMA_signal_248, L8}), .b ({new_AGEMA_signal_264, L10}), .c ({new_AGEMA_signal_276, L27}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L28_U1 ( .a ({new_AGEMA_signal_265, L11}), .b ({new_AGEMA_signal_256, L14}), .c ({new_AGEMA_signal_277, L28}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_L29_U1 ( .a ({new_AGEMA_signal_265, L11}), .b ({new_AGEMA_signal_258, L17}), .c ({new_AGEMA_signal_278, L29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S0_U1 ( .a ({new_AGEMA_signal_261, L6}), .b ({new_AGEMA_signal_273, L24}), .c ({new_AGEMA_signal_280, O[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S1_U1 ( .a ({new_AGEMA_signal_270, L16}), .b ({new_AGEMA_signal_275, L26}), .c ({new_AGEMA_signal_281, O[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S2_U1 ( .a ({new_AGEMA_signal_266, L19}), .b ({new_AGEMA_signal_277, L28}), .c ({new_AGEMA_signal_282, O[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S3_U1 ( .a ({new_AGEMA_signal_261, L6}), .b ({new_AGEMA_signal_272, L21}), .c ({new_AGEMA_signal_283, O[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S4_U1 ( .a ({new_AGEMA_signal_271, L20}), .b ({new_AGEMA_signal_267, L22}), .c ({new_AGEMA_signal_284, O[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S5_U1 ( .a ({new_AGEMA_signal_274, L25}), .b ({new_AGEMA_signal_278, L29}), .c ({new_AGEMA_signal_285, O[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S6_U1 ( .a ({new_AGEMA_signal_269, L13}), .b ({new_AGEMA_signal_276, L27}), .c ({new_AGEMA_signal_286, O[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) XOR_S7_U1 ( .a ({new_AGEMA_signal_261, L6}), .b ({new_AGEMA_signal_268, L23}), .c ({new_AGEMA_signal_279, O[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_7_ ( .clk (clk), .D ({new_AGEMA_signal_280, O[7]}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_6_ ( .clk (clk), .D ({new_AGEMA_signal_281, O[6]}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_5_ ( .clk (clk), .D ({new_AGEMA_signal_282, O[5]}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_4_ ( .clk (clk), .D ({new_AGEMA_signal_283, O[4]}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_3_ ( .clk (clk), .D ({new_AGEMA_signal_284, O[3]}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_2_ ( .clk (clk), .D ({new_AGEMA_signal_285, O[2]}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_1_ ( .clk (clk), .D ({new_AGEMA_signal_286, O[1]}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) Y_reg_0_ ( .clk (clk), .D ({new_AGEMA_signal_279, O[0]}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
