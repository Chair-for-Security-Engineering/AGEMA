
module sbox ( SI, clk, SO );
  (* AGEMA = "secure" *) input [7:0] SI;
  (* AGEMA = "clock" *)  input clk;

  output [7:0] SO;

  wire   N169, N277, N379, N470, N563, N639, N723, N789, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832;

  DFF_X1 SO_reg_7_ ( .D(N169), .CK(clk), .Q(SO[7]), .QN() );
  DFF_X1 SO_reg_6_ ( .D(N277), .CK(clk), .Q(SO[6]), .QN() );
  DFF_X1 SO_reg_5_ ( .D(N379), .CK(clk), .Q(SO[5]), .QN() );
  DFF_X1 SO_reg_4_ ( .D(N470), .CK(clk), .Q(SO[4]), .QN() );
  DFF_X1 SO_reg_3_ ( .D(N563), .CK(clk), .Q(SO[3]), .QN() );
  DFF_X1 SO_reg_2_ ( .D(N639), .CK(clk), .Q(SO[2]), .QN() );
  DFF_X1 SO_reg_1_ ( .D(N723), .CK(clk), .Q(SO[1]), .QN() );
  DFF_X1 SO_reg_0_ ( .D(N789), .CK(clk), .Q(SO[0]), .QN() );
  NOR2_X2 U1937 ( .A1(n2796), .A2(SI[6]), .ZN(n2719) );
  INV_X1 U1938 ( .A(SI[7]), .ZN(n2796) );
  INV_X1 U1939 ( .A(SI[5]), .ZN(n2810) );
  INV_X1 U1940 ( .A(SI[6]), .ZN(n2462) );
  INV_X1 U1941 ( .A(SI[3]), .ZN(n2760) );
  INV_X1 U1942 ( .A(SI[4]), .ZN(n2791) );
  INV_X1 U1943 ( .A(n2624), .ZN(n2672) );
  INV_X1 U1944 ( .A(SI[1]), .ZN(n2813) );
  INV_X1 U1945 ( .A(SI[0]), .ZN(n2630) );
  INV_X1 U1946 ( .A(SI[2]), .ZN(n2765) );
  NAND2_X1 U1947 ( .A1(SI[2]), .A2(SI[3]), .ZN(n2635) );
  NOR2_X1 U1948 ( .A1(n2462), .A2(SI[7]), .ZN(n2641) );
  NOR2_X1 U1949 ( .A1(SI[6]), .A2(SI[5]), .ZN(n2790) );
  NAND2_X1 U1950 ( .A1(SI[6]), .A2(SI[7]), .ZN(n2519) );
  INV_X1 U1951 ( .A(n2519), .ZN(n2750) );
  NAND2_X1 U1952 ( .A1(n2760), .A2(SI[5]), .ZN(n2615) );
  INV_X1 U1953 ( .A(n2615), .ZN(n2640) );
  NAND2_X1 U1954 ( .A1(n2750), .A2(n2640), .ZN(n2575) );
  NAND2_X1 U1955 ( .A1(n2765), .A2(n2630), .ZN(n2699) );
  INV_X1 U1956 ( .A(n2699), .ZN(n2737) );
  NAND2_X1 U1957 ( .A1(n2765), .A2(n2813), .ZN(n2816) );
  INV_X1 U1958 ( .A(n2816), .ZN(n2767) );
  NOR2_X1 U1959 ( .A1(n2737), .A2(n2767), .ZN(n1962) );
  NOR2_X1 U1960 ( .A1(n2575), .A2(n1962), .ZN(n1924) );
  NAND2_X1 U1961 ( .A1(n2765), .A2(SI[1]), .ZN(n2780) );
  INV_X1 U1962 ( .A(n2780), .ZN(n2789) );
  NOR2_X1 U1963 ( .A1(SI[6]), .A2(n2810), .ZN(n2317) );
  NAND2_X1 U1964 ( .A1(n2789), .A2(n2317), .ZN(n1922) );
  NOR2_X1 U1965 ( .A1(n2791), .A2(n2760), .ZN(n2694) );
  INV_X1 U1966 ( .A(n2694), .ZN(n2769) );
  NOR2_X1 U1967 ( .A1(n1922), .A2(n2769), .ZN(n1923) );
  NOR2_X1 U1968 ( .A1(n1924), .A2(n1923), .ZN(n1936) );
  NOR2_X1 U1969 ( .A1(n2760), .A2(SI[4]), .ZN(n2073) );
  INV_X1 U1970 ( .A(n2073), .ZN(n2707) );
  NAND2_X1 U1971 ( .A1(SI[7]), .A2(SI[5]), .ZN(n2315) );
  NOR2_X1 U1972 ( .A1(SI[0]), .A2(SI[1]), .ZN(n2682) );
  INV_X1 U1973 ( .A(n2682), .ZN(n2713) );
  NOR2_X1 U1974 ( .A1(n2315), .A2(n2713), .ZN(n2755) );
  NAND2_X1 U1975 ( .A1(n2813), .A2(SI[0]), .ZN(n2723) );
  INV_X1 U1976 ( .A(n2723), .ZN(n2688) );
  NAND2_X1 U1977 ( .A1(n2317), .A2(n2688), .ZN(n1926) );
  NAND2_X1 U1978 ( .A1(n2810), .A2(SI[7]), .ZN(n2725) );
  INV_X1 U1979 ( .A(n2725), .ZN(n2541) );
  NAND2_X1 U1980 ( .A1(n2767), .A2(n2541), .ZN(n1925) );
  NAND2_X1 U1981 ( .A1(n1926), .A2(n1925), .ZN(n1927) );
  NOR2_X1 U1982 ( .A1(n2755), .A2(n1927), .ZN(n1928) );
  NOR2_X1 U1983 ( .A1(n2707), .A2(n1928), .ZN(n1934) );
  NAND2_X1 U1984 ( .A1(n2760), .A2(SI[4]), .ZN(n2815) );
  INV_X1 U1985 ( .A(n2815), .ZN(n2086) );
  NAND2_X1 U1986 ( .A1(n2086), .A2(n2317), .ZN(n2151) );
  NOR2_X1 U1987 ( .A1(n2810), .A2(n2791), .ZN(n2600) );
  NAND2_X1 U1988 ( .A1(n2641), .A2(n2600), .ZN(n2631) );
  INV_X1 U1989 ( .A(n2631), .ZN(n2734) );
  NOR2_X1 U1990 ( .A1(n2462), .A2(SI[5]), .ZN(n2538) );
  INV_X1 U1991 ( .A(n2538), .ZN(n2786) );
  NOR2_X1 U1992 ( .A1(n2707), .A2(n2786), .ZN(n2763) );
  NOR2_X1 U1993 ( .A1(n2734), .A2(n2763), .ZN(n1929) );
  NAND2_X1 U1994 ( .A1(n2151), .A2(n1929), .ZN(n1931) );
  NOR2_X1 U1995 ( .A1(SI[4]), .A2(SI[3]), .ZN(n2595) );
  INV_X1 U1996 ( .A(n2595), .ZN(n2742) );
  NOR2_X1 U1997 ( .A1(n2519), .A2(n2742), .ZN(n1930) );
  NOR2_X1 U1998 ( .A1(n1931), .A2(n1930), .ZN(n1932) );
  NOR2_X1 U1999 ( .A1(n2765), .A2(n2630), .ZN(n2753) );
  INV_X1 U2000 ( .A(n2753), .ZN(n2577) );
  NOR2_X1 U2001 ( .A1(n1932), .A2(n2577), .ZN(n1933) );
  NOR2_X1 U2002 ( .A1(n1934), .A2(n1933), .ZN(n1935) );
  NAND2_X1 U2003 ( .A1(n1936), .A2(n1935), .ZN(n1941) );
  NAND2_X1 U2004 ( .A1(n2810), .A2(SI[4]), .ZN(n2400) );
  NOR2_X1 U2005 ( .A1(n2400), .A2(n2519), .ZN(n2492) );
  INV_X1 U2006 ( .A(n2492), .ZN(n2732) );
  NOR2_X1 U2007 ( .A1(SI[3]), .A2(n2732), .ZN(n2665) );
  NAND2_X1 U2008 ( .A1(n2765), .A2(SI[3]), .ZN(n2785) );
  INV_X1 U2009 ( .A(n2785), .ZN(n2792) );
  NAND2_X1 U2010 ( .A1(SI[4]), .A2(n2792), .ZN(n1937) );
  NOR2_X1 U2011 ( .A1(SI[6]), .A2(n1937), .ZN(n1938) );
  NOR2_X1 U2012 ( .A1(n2665), .A2(n1938), .ZN(n1939) );
  NOR2_X1 U2013 ( .A1(n2813), .A2(SI[0]), .ZN(n2609) );
  INV_X1 U2014 ( .A(n2609), .ZN(n2724) );
  NOR2_X1 U2015 ( .A1(n1939), .A2(n2724), .ZN(n1940) );
  NOR2_X1 U2016 ( .A1(n1941), .A2(n1940), .ZN(n2019) );
  NOR2_X1 U2017 ( .A1(n2760), .A2(n2813), .ZN(n2661) );
  INV_X1 U2018 ( .A(n2661), .ZN(n2174) );
  NOR2_X1 U2019 ( .A1(n2174), .A2(n2732), .ZN(n2235) );
  NAND2_X1 U2020 ( .A1(SI[2]), .A2(SI[1]), .ZN(n2708) );
  INV_X1 U2021 ( .A(n2708), .ZN(n2493) );
  NAND2_X1 U2022 ( .A1(SI[6]), .A2(n2493), .ZN(n1942) );
  NOR2_X1 U2023 ( .A1(SI[4]), .A2(n1942), .ZN(n1943) );
  NOR2_X1 U2024 ( .A1(n2235), .A2(n1943), .ZN(n1948) );
  NAND2_X1 U2025 ( .A1(n2796), .A2(SI[5]), .ZN(n2587) );
  OR2_X1 U2026 ( .A1(n2587), .A2(n2815), .ZN(n2676) );
  NAND2_X1 U2027 ( .A1(n2676), .A2(SI[0]), .ZN(n1946) );
  INV_X1 U2028 ( .A(n2719), .ZN(n2570) );
  NOR2_X1 U2029 ( .A1(SI[5]), .A2(SI[3]), .ZN(n2559) );
  NAND2_X1 U2030 ( .A1(n2789), .A2(n2559), .ZN(n1944) );
  NOR2_X1 U2031 ( .A1(n2570), .A2(n1944), .ZN(n1945) );
  NOR2_X1 U2032 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
  NAND2_X1 U2033 ( .A1(n1948), .A2(n1947), .ZN(n1961) );
  NAND2_X1 U2034 ( .A1(n2792), .A2(n2734), .ZN(n1956) );
  NOR2_X1 U2035 ( .A1(n2765), .A2(SI[1]), .ZN(n2643) );
  INV_X1 U2036 ( .A(n2643), .ZN(n2442) );
  NOR2_X1 U2037 ( .A1(n2725), .A2(n2769), .ZN(n1950) );
  INV_X1 U2038 ( .A(n2790), .ZN(n2739) );
  NOR2_X1 U2039 ( .A1(SI[7]), .A2(n2739), .ZN(n1949) );
  NOR2_X1 U2040 ( .A1(n1950), .A2(n1949), .ZN(n1951) );
  NOR2_X1 U2041 ( .A1(n2442), .A2(n1951), .ZN(n1954) );
  NAND2_X1 U2042 ( .A1(n2750), .A2(n2600), .ZN(n2677) );
  INV_X1 U2043 ( .A(n2677), .ZN(n2662) );
  NAND2_X1 U2044 ( .A1(n2462), .A2(n2796), .ZN(n2437) );
  NOR2_X1 U2045 ( .A1(SI[5]), .A2(SI[4]), .ZN(n2261) );
  INV_X1 U2046 ( .A(n2261), .ZN(n2778) );
  NOR2_X1 U2047 ( .A1(n2437), .A2(n2778), .ZN(n2627) );
  NOR2_X1 U2048 ( .A1(n2662), .A2(n2627), .ZN(n1952) );
  NOR2_X1 U2049 ( .A1(n2635), .A2(n1952), .ZN(n1953) );
  NOR2_X1 U2050 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  NAND2_X1 U2051 ( .A1(n1956), .A2(n1955), .ZN(n1958) );
  NAND2_X1 U2052 ( .A1(SI[7]), .A2(n2791), .ZN(n2452) );
  NOR2_X1 U2053 ( .A1(n2816), .A2(n2452), .ZN(n1957) );
  NOR2_X1 U2054 ( .A1(n1958), .A2(n1957), .ZN(n1959) );
  INV_X1 U2055 ( .A(n2437), .ZN(n2766) );
  NAND2_X1 U2056 ( .A1(n2766), .A2(n2600), .ZN(n2088) );
  NOR2_X1 U2057 ( .A1(n2635), .A2(n2088), .ZN(n2687) );
  NOR2_X1 U2058 ( .A1(SI[0]), .A2(n2687), .ZN(n2658) );
  NAND2_X1 U2059 ( .A1(n1959), .A2(n2658), .ZN(n1960) );
  NAND2_X1 U2060 ( .A1(n1961), .A2(n1960), .ZN(n2002) );
  OR2_X1 U2061 ( .A1(n1962), .A2(n2587), .ZN(n1966) );
  NOR2_X1 U2062 ( .A1(n2519), .A2(n2708), .ZN(n1964) );
  NAND2_X1 U2063 ( .A1(SI[0]), .A2(n2643), .ZN(n2736) );
  NOR2_X1 U2064 ( .A1(n2736), .A2(n2725), .ZN(n1963) );
  NOR2_X1 U2065 ( .A1(n1964), .A2(n1963), .ZN(n1965) );
  NAND2_X1 U2066 ( .A1(n1966), .A2(n1965), .ZN(n1967) );
  NAND2_X1 U2067 ( .A1(n1967), .A2(n2595), .ZN(n1990) );
  NOR2_X1 U2068 ( .A1(n2765), .A2(SI[3]), .ZN(n2772) );
  NAND2_X1 U2069 ( .A1(n2772), .A2(SI[1]), .ZN(n2673) );
  NAND2_X1 U2070 ( .A1(n2791), .A2(SI[5]), .ZN(n2824) );
  INV_X1 U2071 ( .A(n2824), .ZN(n2612) );
  NAND2_X1 U2072 ( .A1(n2766), .A2(n2612), .ZN(n2761) );
  INV_X1 U2073 ( .A(n2761), .ZN(n2720) );
  INV_X1 U2074 ( .A(n2400), .ZN(n2313) );
  NAND2_X1 U2075 ( .A1(n2313), .A2(n2719), .ZN(n2412) );
  INV_X1 U2076 ( .A(n2412), .ZN(n2417) );
  NOR2_X1 U2077 ( .A1(n2720), .A2(n2417), .ZN(n1968) );
  NOR2_X1 U2078 ( .A1(n2673), .A2(n1968), .ZN(n1970) );
  NAND2_X1 U2079 ( .A1(n2641), .A2(n2261), .ZN(n2571) );
  INV_X1 U2080 ( .A(n2571), .ZN(n2505) );
  NOR2_X1 U2081 ( .A1(n2519), .A2(n2824), .ZN(n2651) );
  NOR2_X1 U2082 ( .A1(n2505), .A2(n2651), .ZN(n2684) );
  NAND2_X1 U2083 ( .A1(n2792), .A2(SI[1]), .ZN(n2359) );
  NOR2_X1 U2084 ( .A1(n2684), .A2(n2359), .ZN(n1969) );
  NOR2_X1 U2085 ( .A1(n1970), .A2(n1969), .ZN(n1984) );
  NOR2_X1 U2086 ( .A1(n2519), .A2(n2778), .ZN(n2101) );
  INV_X1 U2087 ( .A(n2101), .ZN(n2625) );
  NOR2_X1 U2088 ( .A1(n2708), .A2(n2625), .ZN(n1972) );
  NOR2_X1 U2089 ( .A1(n2810), .A2(n2760), .ZN(n2395) );
  INV_X1 U2090 ( .A(n2395), .ZN(n2818) );
  NAND2_X1 U2091 ( .A1(n2719), .A2(n2609), .ZN(n2190) );
  NOR2_X1 U2092 ( .A1(n2818), .A2(n2190), .ZN(n1971) );
  NOR2_X1 U2093 ( .A1(n1972), .A2(n1971), .ZN(n1978) );
  NAND2_X1 U2094 ( .A1(SI[6]), .A2(SI[5]), .ZN(n2779) );
  NAND2_X1 U2095 ( .A1(n2739), .A2(n2779), .ZN(n1976) );
  NOR2_X1 U2096 ( .A1(n2630), .A2(n2813), .ZN(n2624) );
  NAND2_X1 U2097 ( .A1(SI[4]), .A2(SI[2]), .ZN(n2242) );
  NOR2_X1 U2098 ( .A1(n2672), .A2(n2242), .ZN(n2535) );
  NAND2_X1 U2099 ( .A1(n2790), .A2(n2535), .ZN(n1974) );
  NOR2_X1 U2100 ( .A1(SI[2]), .A2(n2791), .ZN(n2356) );
  NAND2_X1 U2101 ( .A1(n2688), .A2(n2356), .ZN(n1973) );
  NAND2_X1 U2102 ( .A1(n1974), .A2(n1973), .ZN(n1975) );
  NAND2_X1 U2103 ( .A1(n1976), .A2(n1975), .ZN(n1977) );
  NAND2_X1 U2104 ( .A1(n1978), .A2(n1977), .ZN(n1982) );
  NOR2_X1 U2105 ( .A1(n2815), .A2(n2315), .ZN(n2690) );
  NOR2_X1 U2106 ( .A1(n2732), .A2(n2635), .ZN(n1979) );
  NOR2_X1 U2107 ( .A1(n2690), .A2(n1979), .ZN(n1980) );
  NOR2_X1 U2108 ( .A1(SI[1]), .A2(n1980), .ZN(n1981) );
  NOR2_X1 U2109 ( .A1(n1982), .A2(n1981), .ZN(n1983) );
  NAND2_X1 U2110 ( .A1(n1984), .A2(n1983), .ZN(n1988) );
  NAND2_X1 U2111 ( .A1(n2493), .A2(n2630), .ZN(n2817) );
  NOR2_X1 U2112 ( .A1(n2786), .A2(n2817), .ZN(n1985) );
  NOR2_X1 U2113 ( .A1(n2442), .A2(n2779), .ZN(n2741) );
  NOR2_X1 U2114 ( .A1(n1985), .A2(n2741), .ZN(n1986) );
  NOR2_X1 U2115 ( .A1(n2815), .A2(n1986), .ZN(n1987) );
  NOR2_X1 U2116 ( .A1(n1988), .A2(n1987), .ZN(n1989) );
  NAND2_X1 U2117 ( .A1(n1990), .A2(n1989), .ZN(n2000) );
  NOR2_X1 U2118 ( .A1(n2780), .A2(n2818), .ZN(n1992) );
  INV_X1 U2119 ( .A(n2772), .ZN(n2823) );
  NOR2_X1 U2120 ( .A1(n2823), .A2(n2672), .ZN(n1991) );
  NOR2_X1 U2121 ( .A1(n1992), .A2(n1991), .ZN(n1994) );
  NOR2_X1 U2122 ( .A1(n2760), .A2(SI[5]), .ZN(n2611) );
  NAND2_X1 U2123 ( .A1(n2643), .A2(n2611), .ZN(n1993) );
  NAND2_X1 U2124 ( .A1(n1994), .A2(n1993), .ZN(n1997) );
  NOR2_X1 U2125 ( .A1(n2737), .A2(n2792), .ZN(n1995) );
  NOR2_X1 U2126 ( .A1(n2400), .A2(n1995), .ZN(n1996) );
  NOR2_X1 U2127 ( .A1(n1997), .A2(n1996), .ZN(n1998) );
  NOR2_X1 U2128 ( .A1(n2437), .A2(n1998), .ZN(n1999) );
  NOR2_X1 U2129 ( .A1(n2000), .A2(n1999), .ZN(n2001) );
  NAND2_X1 U2130 ( .A1(n2002), .A2(n2001), .ZN(n2017) );
  INV_X1 U2131 ( .A(n2641), .ZN(n2828) );
  NOR2_X1 U2132 ( .A1(n2818), .A2(n2708), .ZN(n2241) );
  NAND2_X1 U2133 ( .A1(n2765), .A2(SI[0]), .ZN(n2616) );
  INV_X1 U2134 ( .A(n2616), .ZN(n2679) );
  NAND2_X1 U2135 ( .A1(SI[5]), .A2(n2679), .ZN(n2003) );
  NOR2_X1 U2136 ( .A1(SI[1]), .A2(n2003), .ZN(n2137) );
  NOR2_X1 U2137 ( .A1(n2241), .A2(n2137), .ZN(n2012) );
  NAND2_X1 U2138 ( .A1(n2765), .A2(n2760), .ZN(n2563) );
  INV_X1 U2139 ( .A(n2563), .ZN(n2809) );
  NAND2_X1 U2140 ( .A1(n2612), .A2(n2809), .ZN(n2008) );
  NOR2_X1 U2141 ( .A1(n2679), .A2(n2688), .ZN(n2572) );
  NOR2_X1 U2142 ( .A1(n2815), .A2(n2572), .ZN(n2006) );
  NOR2_X1 U2143 ( .A1(n2809), .A2(n2356), .ZN(n2004) );
  NOR2_X1 U2144 ( .A1(n2723), .A2(n2004), .ZN(n2005) );
  NOR2_X1 U2145 ( .A1(n2006), .A2(n2005), .ZN(n2007) );
  NAND2_X1 U2146 ( .A1(n2008), .A2(n2007), .ZN(n2010) );
  NOR2_X1 U2147 ( .A1(n2635), .A2(n2672), .ZN(n2009) );
  NOR2_X1 U2148 ( .A1(n2010), .A2(n2009), .ZN(n2011) );
  NAND2_X1 U2149 ( .A1(n2012), .A2(n2011), .ZN(n2014) );
  INV_X1 U2150 ( .A(n2611), .ZN(n2709) );
  NAND2_X1 U2151 ( .A1(n2789), .A2(n2630), .ZN(n2533) );
  NOR2_X1 U2152 ( .A1(n2709), .A2(n2533), .ZN(n2013) );
  NOR2_X1 U2153 ( .A1(n2014), .A2(n2013), .ZN(n2015) );
  NOR2_X1 U2154 ( .A1(n2828), .A2(n2015), .ZN(n2016) );
  NOR2_X1 U2155 ( .A1(n2017), .A2(n2016), .ZN(n2018) );
  NAND2_X1 U2156 ( .A1(n2019), .A2(n2018), .ZN(N169) );
  NAND2_X1 U2157 ( .A1(n2719), .A2(n2682), .ZN(n2026) );
  NAND2_X1 U2158 ( .A1(n2766), .A2(n2493), .ZN(n2022) );
  NOR2_X1 U2159 ( .A1(n2462), .A2(n2725), .ZN(n2227) );
  NAND2_X1 U2160 ( .A1(n2753), .A2(n2227), .ZN(n2020) );
  MUX2_X1 U2161 ( .A(n2020), .B(n2779), .S(n2813), .Z(n2021) );
  NAND2_X1 U2162 ( .A1(n2022), .A2(n2021), .ZN(n2024) );
  NAND2_X1 U2163 ( .A1(n2796), .A2(n2810), .ZN(n2401) );
  NOR2_X1 U2164 ( .A1(n2817), .A2(n2401), .ZN(n2023) );
  NOR2_X1 U2165 ( .A1(n2024), .A2(n2023), .ZN(n2025) );
  NAND2_X1 U2166 ( .A1(n2026), .A2(n2025), .ZN(n2029) );
  NAND2_X1 U2167 ( .A1(n2790), .A2(n2630), .ZN(n2027) );
  NOR2_X1 U2168 ( .A1(n2027), .A2(n2765), .ZN(n2028) );
  NOR2_X1 U2169 ( .A1(n2029), .A2(n2028), .ZN(n2030) );
  NOR2_X1 U2170 ( .A1(n2742), .A2(n2030), .ZN(n2038) );
  NOR2_X1 U2171 ( .A1(n2818), .A2(n2442), .ZN(n2214) );
  NAND2_X1 U2172 ( .A1(n2214), .A2(n2630), .ZN(n2033) );
  NOR2_X1 U2173 ( .A1(n2442), .A2(n2707), .ZN(n2290) );
  NAND2_X1 U2174 ( .A1(SI[0]), .A2(n2767), .ZN(n2376) );
  NOR2_X1 U2175 ( .A1(n2376), .A2(n2615), .ZN(n2031) );
  NOR2_X1 U2176 ( .A1(n2290), .A2(n2031), .ZN(n2032) );
  NAND2_X1 U2177 ( .A1(n2033), .A2(n2032), .ZN(n2035) );
  NOR2_X1 U2178 ( .A1(n2708), .A2(n2400), .ZN(n2034) );
  NOR2_X1 U2179 ( .A1(n2035), .A2(n2034), .ZN(n2036) );
  NOR2_X1 U2180 ( .A1(n2437), .A2(n2036), .ZN(n2037) );
  NOR2_X1 U2181 ( .A1(n2038), .A2(n2037), .ZN(n2113) );
  NAND2_X1 U2182 ( .A1(n2611), .A2(n2719), .ZN(n2171) );
  NOR2_X1 U2183 ( .A1(n2828), .A2(n2769), .ZN(n2039) );
  NOR2_X1 U2184 ( .A1(n2627), .A2(n2039), .ZN(n2040) );
  NAND2_X1 U2185 ( .A1(n2171), .A2(n2040), .ZN(n2041) );
  NAND2_X1 U2186 ( .A1(n2041), .A2(n2753), .ZN(n2054) );
  NAND2_X1 U2187 ( .A1(n2643), .A2(n2651), .ZN(n2050) );
  NOR2_X1 U2188 ( .A1(n2725), .A2(n2707), .ZN(n2042) );
  NOR2_X1 U2189 ( .A1(n2665), .A2(n2042), .ZN(n2043) );
  NOR2_X1 U2190 ( .A1(n2713), .A2(n2043), .ZN(n2048) );
  NOR2_X1 U2191 ( .A1(n2707), .A2(n2315), .ZN(n2754) );
  NOR2_X1 U2192 ( .A1(n2313), .A2(n2790), .ZN(n2044) );
  NOR2_X1 U2193 ( .A1(n2563), .A2(n2044), .ZN(n2045) );
  NOR2_X1 U2194 ( .A1(n2754), .A2(n2045), .ZN(n2046) );
  NOR2_X1 U2195 ( .A1(n2046), .A2(n2672), .ZN(n2047) );
  NOR2_X1 U2196 ( .A1(n2048), .A2(n2047), .ZN(n2049) );
  NAND2_X1 U2197 ( .A1(n2050), .A2(n2049), .ZN(n2052) );
  NAND2_X1 U2198 ( .A1(n2313), .A2(n2641), .ZN(n2654) );
  NOR2_X1 U2199 ( .A1(n2654), .A2(n2635), .ZN(n2051) );
  NOR2_X1 U2200 ( .A1(n2052), .A2(n2051), .ZN(n2053) );
  NAND2_X1 U2201 ( .A1(n2054), .A2(n2053), .ZN(n2111) );
  NAND2_X1 U2202 ( .A1(n2635), .A2(n2577), .ZN(n2055) );
  NAND2_X1 U2203 ( .A1(n2612), .A2(n2055), .ZN(n2056) );
  MUX2_X1 U2204 ( .A(n2056), .B(n2769), .S(n2813), .Z(n2058) );
  NAND2_X1 U2205 ( .A1(n2395), .A2(n2767), .ZN(n2057) );
  NAND2_X1 U2206 ( .A1(n2058), .A2(n2057), .ZN(n2059) );
  NAND2_X1 U2207 ( .A1(n2719), .A2(n2059), .ZN(n2072) );
  NOR2_X1 U2208 ( .A1(n2679), .A2(n2682), .ZN(n2407) );
  NOR2_X1 U2209 ( .A1(n2407), .A2(n2824), .ZN(n2060) );
  NOR2_X1 U2210 ( .A1(n2535), .A2(n2060), .ZN(n2063) );
  NOR2_X1 U2211 ( .A1(n2765), .A2(SI[5]), .ZN(n2061) );
  NAND2_X1 U2212 ( .A1(n2688), .A2(n2061), .ZN(n2062) );
  NAND2_X1 U2213 ( .A1(n2063), .A2(n2062), .ZN(n2064) );
  NAND2_X1 U2214 ( .A1(n2641), .A2(n2064), .ZN(n2067) );
  NOR2_X1 U2215 ( .A1(n2816), .A2(n2654), .ZN(n2066) );
  NAND2_X1 U2216 ( .A1(n2766), .A2(n2559), .ZN(n2731) );
  NOR2_X1 U2217 ( .A1(n2765), .A2(n2731), .ZN(n2065) );
  NOR2_X1 U2218 ( .A1(n2066), .A2(n2065), .ZN(n2652) );
  NAND2_X1 U2219 ( .A1(n2067), .A2(n2652), .ZN(n2070) );
  INV_X1 U2220 ( .A(n2690), .ZN(n2068) );
  NOR2_X1 U2221 ( .A1(n2068), .A2(n2817), .ZN(n2069) );
  NOR2_X1 U2222 ( .A1(n2070), .A2(n2069), .ZN(n2071) );
  NAND2_X1 U2223 ( .A1(n2072), .A2(n2071), .ZN(n2079) );
  NAND2_X1 U2224 ( .A1(n2611), .A2(n2750), .ZN(n2642) );
  NAND2_X1 U2225 ( .A1(n2725), .A2(n2786), .ZN(n2252) );
  NAND2_X1 U2226 ( .A1(n2073), .A2(n2252), .ZN(n2074) );
  NAND2_X1 U2227 ( .A1(n2642), .A2(n2074), .ZN(n2076) );
  NOR2_X1 U2228 ( .A1(n2739), .A2(n2815), .ZN(n2075) );
  NOR2_X1 U2229 ( .A1(n2076), .A2(n2075), .ZN(n2077) );
  NOR2_X1 U2230 ( .A1(n2699), .A2(n2077), .ZN(n2078) );
  NOR2_X1 U2231 ( .A1(n2079), .A2(n2078), .ZN(n2109) );
  NOR2_X1 U2232 ( .A1(n2796), .A2(n2791), .ZN(n2721) );
  OR2_X1 U2233 ( .A1(n2635), .A2(n2723), .ZN(n2081) );
  NAND2_X1 U2234 ( .A1(n2792), .A2(n2682), .ZN(n2080) );
  NAND2_X1 U2235 ( .A1(n2081), .A2(n2080), .ZN(n2082) );
  NAND2_X1 U2236 ( .A1(n2721), .A2(n2082), .ZN(n2105) );
  NAND2_X1 U2237 ( .A1(n2600), .A2(n2719), .ZN(n2498) );
  INV_X1 U2238 ( .A(n2498), .ZN(n2773) );
  NOR2_X1 U2239 ( .A1(n2767), .A2(n2792), .ZN(n2083) );
  NAND2_X1 U2240 ( .A1(n2723), .A2(n2083), .ZN(n2084) );
  NAND2_X1 U2241 ( .A1(n2773), .A2(n2084), .ZN(n2099) );
  NAND2_X1 U2242 ( .A1(n2533), .A2(SI[3]), .ZN(n2085) );
  NAND2_X1 U2243 ( .A1(n2085), .A2(n2627), .ZN(n2091) );
  NAND2_X1 U2244 ( .A1(SI[5]), .A2(n2086), .ZN(n2562) );
  NOR2_X1 U2245 ( .A1(n2519), .A2(n2562), .ZN(n2131) );
  AND2_X1 U2246 ( .A1(n2753), .A2(n2131), .ZN(n2090) );
  NAND2_X1 U2247 ( .A1(SI[0]), .A2(n2661), .ZN(n2087) );
  NOR2_X1 U2248 ( .A1(n2088), .A2(n2087), .ZN(n2089) );
  NOR2_X1 U2249 ( .A1(n2090), .A2(n2089), .ZN(n2158) );
  NAND2_X1 U2250 ( .A1(n2091), .A2(n2158), .ZN(n2097) );
  NAND2_X1 U2251 ( .A1(n2563), .A2(n2174), .ZN(n2156) );
  NAND2_X1 U2252 ( .A1(n2630), .A2(n2156), .ZN(n2330) );
  NOR2_X1 U2253 ( .A1(n2631), .A2(n2330), .ZN(n2093) );
  NOR2_X1 U2254 ( .A1(n2616), .A2(n2151), .ZN(n2092) );
  NOR2_X1 U2255 ( .A1(n2093), .A2(n2092), .ZN(n2095) );
  OR2_X1 U2256 ( .A1(n2761), .A2(n2359), .ZN(n2094) );
  NAND2_X1 U2257 ( .A1(n2095), .A2(n2094), .ZN(n2096) );
  NOR2_X1 U2258 ( .A1(n2097), .A2(n2096), .ZN(n2098) );
  NAND2_X1 U2259 ( .A1(n2099), .A2(n2098), .ZN(n2103) );
  NOR2_X1 U2260 ( .A1(n2769), .A2(n2401), .ZN(n2100) );
  NOR2_X1 U2261 ( .A1(n2101), .A2(n2100), .ZN(n2160) );
  NOR2_X1 U2262 ( .A1(n2376), .A2(n2160), .ZN(n2102) );
  NOR2_X1 U2263 ( .A1(n2103), .A2(n2102), .ZN(n2104) );
  NAND2_X1 U2264 ( .A1(n2105), .A2(n2104), .ZN(n2107) );
  NAND2_X1 U2265 ( .A1(n2492), .A2(n2630), .ZN(n2504) );
  NOR2_X1 U2266 ( .A1(n2504), .A2(n2823), .ZN(n2106) );
  NOR2_X1 U2267 ( .A1(n2107), .A2(n2106), .ZN(n2108) );
  NAND2_X1 U2268 ( .A1(n2109), .A2(n2108), .ZN(n2110) );
  NOR2_X1 U2269 ( .A1(n2111), .A2(n2110), .ZN(n2112) );
  NAND2_X1 U2270 ( .A1(n2113), .A2(n2112), .ZN(N277) );
  NOR2_X1 U2271 ( .A1(n2417), .A2(n2651), .ZN(n2114) );
  NOR2_X1 U2272 ( .A1(n2713), .A2(n2114), .ZN(n2116) );
  NOR2_X1 U2273 ( .A1(n2677), .A2(n2723), .ZN(n2115) );
  NOR2_X1 U2274 ( .A1(n2116), .A2(n2115), .ZN(n2117) );
  NOR2_X1 U2275 ( .A1(SI[3]), .A2(n2117), .ZN(n2128) );
  NAND2_X1 U2276 ( .A1(n2791), .A2(n2765), .ZN(n2298) );
  NOR2_X1 U2277 ( .A1(n2739), .A2(n2298), .ZN(n2544) );
  INV_X1 U2278 ( .A(n2401), .ZN(n2118) );
  NAND2_X1 U2279 ( .A1(n2356), .A2(n2118), .ZN(n2121) );
  NOR2_X1 U2280 ( .A1(n2791), .A2(n2731), .ZN(n2291) );
  NOR2_X1 U2281 ( .A1(SI[3]), .A2(n2498), .ZN(n2119) );
  NOR2_X1 U2282 ( .A1(n2291), .A2(n2119), .ZN(n2120) );
  NAND2_X1 U2283 ( .A1(n2121), .A2(n2120), .ZN(n2123) );
  NOR2_X1 U2284 ( .A1(n2707), .A2(n2570), .ZN(n2122) );
  NOR2_X1 U2285 ( .A1(n2123), .A2(n2122), .ZN(n2124) );
  NAND2_X1 U2286 ( .A1(n2792), .A2(n2612), .ZN(n2811) );
  NAND2_X1 U2287 ( .A1(n2124), .A2(n2811), .ZN(n2125) );
  NOR2_X1 U2288 ( .A1(n2544), .A2(n2125), .ZN(n2126) );
  NOR2_X1 U2289 ( .A1(n2672), .A2(n2126), .ZN(n2127) );
  NOR2_X1 U2290 ( .A1(n2128), .A2(n2127), .ZN(n2212) );
  NOR2_X1 U2291 ( .A1(n2780), .A2(n2498), .ZN(n2130) );
  NOR2_X1 U2292 ( .A1(n2817), .A2(n2631), .ZN(n2129) );
  NOR2_X1 U2293 ( .A1(n2130), .A2(n2129), .ZN(n2155) );
  NOR2_X1 U2294 ( .A1(n2437), .A2(n2742), .ZN(n2647) );
  NAND2_X1 U2295 ( .A1(n2647), .A2(n2813), .ZN(n2150) );
  NAND2_X1 U2296 ( .A1(n2643), .A2(n2131), .ZN(n2543) );
  NOR2_X1 U2297 ( .A1(n2742), .A2(n2315), .ZN(n2132) );
  NOR2_X1 U2298 ( .A1(n2492), .A2(n2132), .ZN(n2133) );
  NOR2_X1 U2299 ( .A1(n2133), .A2(n2816), .ZN(n2134) );
  NOR2_X1 U2300 ( .A1(n2687), .A2(n2134), .ZN(n2135) );
  NAND2_X1 U2301 ( .A1(n2543), .A2(n2135), .ZN(n2148) );
  NOR2_X1 U2302 ( .A1(n2533), .A2(n2742), .ZN(n2136) );
  NOR2_X1 U2303 ( .A1(n2137), .A2(n2136), .ZN(n2143) );
  NOR2_X1 U2304 ( .A1(n2616), .A2(n2707), .ZN(n2220) );
  NAND2_X1 U2305 ( .A1(SI[4]), .A2(n2767), .ZN(n2138) );
  NAND2_X1 U2306 ( .A1(n2572), .A2(n2138), .ZN(n2139) );
  NOR2_X1 U2307 ( .A1(SI[4]), .A2(n2630), .ZN(n2346) );
  NOR2_X1 U2308 ( .A1(n2139), .A2(n2346), .ZN(n2140) );
  NOR2_X1 U2309 ( .A1(n2818), .A2(n2140), .ZN(n2141) );
  NOR2_X1 U2310 ( .A1(n2220), .A2(n2141), .ZN(n2142) );
  NAND2_X1 U2311 ( .A1(n2143), .A2(n2142), .ZN(n2145) );
  NAND2_X1 U2312 ( .A1(n2612), .A2(n2760), .ZN(n2555) );
  NOR2_X1 U2313 ( .A1(n2724), .A2(n2555), .ZN(n2144) );
  NOR2_X1 U2314 ( .A1(n2145), .A2(n2144), .ZN(n2146) );
  NOR2_X1 U2315 ( .A1(n2828), .A2(n2146), .ZN(n2147) );
  NOR2_X1 U2316 ( .A1(n2148), .A2(n2147), .ZN(n2149) );
  NAND2_X1 U2317 ( .A1(n2150), .A2(n2149), .ZN(n2153) );
  NOR2_X1 U2318 ( .A1(n2151), .A2(n2533), .ZN(n2152) );
  NOR2_X1 U2319 ( .A1(n2153), .A2(n2152), .ZN(n2154) );
  NAND2_X1 U2320 ( .A1(n2155), .A2(n2154), .ZN(n2210) );
  NAND2_X1 U2321 ( .A1(n2627), .A2(n2156), .ZN(n2170) );
  NAND2_X1 U2322 ( .A1(n2612), .A2(n2796), .ZN(n2429) );
  NAND2_X1 U2323 ( .A1(n2429), .A2(n2732), .ZN(n2157) );
  NAND2_X1 U2324 ( .A1(n2157), .A2(n2679), .ZN(n2159) );
  NAND2_X1 U2325 ( .A1(n2159), .A2(n2158), .ZN(n2168) );
  NAND2_X1 U2326 ( .A1(n2160), .A2(n2498), .ZN(n2161) );
  NAND2_X1 U2327 ( .A1(n2737), .A2(n2161), .ZN(n2166) );
  NOR2_X1 U2328 ( .A1(n2437), .A2(n2630), .ZN(n2162) );
  NOR2_X1 U2329 ( .A1(n2317), .A2(n2162), .ZN(n2163) );
  NOR2_X1 U2330 ( .A1(n2442), .A2(n2163), .ZN(n2164) );
  NAND2_X1 U2331 ( .A1(n2694), .A2(n2164), .ZN(n2165) );
  NAND2_X1 U2332 ( .A1(n2166), .A2(n2165), .ZN(n2167) );
  NOR2_X1 U2333 ( .A1(n2168), .A2(n2167), .ZN(n2169) );
  NAND2_X1 U2334 ( .A1(n2170), .A2(n2169), .ZN(n2173) );
  NOR2_X1 U2335 ( .A1(n2171), .A2(n2376), .ZN(n2172) );
  NOR2_X1 U2336 ( .A1(n2173), .A2(n2172), .ZN(n2208) );
  NOR2_X1 U2337 ( .A1(n2315), .A2(n2242), .ZN(n2545) );
  NAND2_X1 U2338 ( .A1(SI[3]), .A2(n2545), .ZN(n2186) );
  NAND2_X1 U2339 ( .A1(n2790), .A2(n2290), .ZN(n2181) );
  NAND2_X1 U2340 ( .A1(n2559), .A2(n2643), .ZN(n2178) );
  NAND2_X1 U2341 ( .A1(SI[2]), .A2(n2791), .ZN(n2430) );
  NAND2_X1 U2342 ( .A1(n2430), .A2(n2707), .ZN(n2176) );
  NOR2_X1 U2343 ( .A1(n2174), .A2(SI[5]), .ZN(n2175) );
  NOR2_X1 U2344 ( .A1(n2176), .A2(n2175), .ZN(n2177) );
  NAND2_X1 U2345 ( .A1(n2178), .A2(n2177), .ZN(n2179) );
  NAND2_X1 U2346 ( .A1(n2179), .A2(n2766), .ZN(n2180) );
  NAND2_X1 U2347 ( .A1(n2181), .A2(n2180), .ZN(n2184) );
  NAND2_X1 U2348 ( .A1(n2261), .A2(n2796), .ZN(n2182) );
  NOR2_X1 U2349 ( .A1(n2635), .A2(n2182), .ZN(n2183) );
  NOR2_X1 U2350 ( .A1(n2184), .A2(n2183), .ZN(n2185) );
  NAND2_X1 U2351 ( .A1(n2186), .A2(n2185), .ZN(n2187) );
  NAND2_X1 U2352 ( .A1(n2187), .A2(n2630), .ZN(n2199) );
  NOR2_X1 U2353 ( .A1(n2786), .A2(n2430), .ZN(n2188) );
  NAND2_X1 U2354 ( .A1(n2688), .A2(n2188), .ZN(n2195) );
  NOR2_X1 U2355 ( .A1(n2792), .A2(n2612), .ZN(n2189) );
  NOR2_X1 U2356 ( .A1(n2190), .A2(n2189), .ZN(n2193) );
  NAND2_X1 U2357 ( .A1(n2635), .A2(n2769), .ZN(n2446) );
  NAND2_X1 U2358 ( .A1(n2609), .A2(n2446), .ZN(n2191) );
  NOR2_X1 U2359 ( .A1(n2315), .A2(n2191), .ZN(n2192) );
  NOR2_X1 U2360 ( .A1(n2193), .A2(n2192), .ZN(n2194) );
  NAND2_X1 U2361 ( .A1(n2195), .A2(n2194), .ZN(n2197) );
  NAND2_X1 U2362 ( .A1(n2750), .A2(n2559), .ZN(n2576) );
  NOR2_X1 U2363 ( .A1(n2609), .A2(n2765), .ZN(n2748) );
  NOR2_X1 U2364 ( .A1(n2576), .A2(n2748), .ZN(n2196) );
  NOR2_X1 U2365 ( .A1(n2197), .A2(n2196), .ZN(n2198) );
  NAND2_X1 U2366 ( .A1(n2199), .A2(n2198), .ZN(n2206) );
  NAND2_X1 U2367 ( .A1(SI[0]), .A2(n2505), .ZN(n2201) );
  INV_X1 U2368 ( .A(n2654), .ZN(n2674) );
  NAND2_X1 U2369 ( .A1(n2674), .A2(n2672), .ZN(n2200) );
  NAND2_X1 U2370 ( .A1(n2201), .A2(n2200), .ZN(n2203) );
  MUX2_X1 U2371 ( .A(n2734), .B(n2417), .S(n2813), .Z(n2202) );
  NOR2_X1 U2372 ( .A1(n2203), .A2(n2202), .ZN(n2204) );
  NOR2_X1 U2373 ( .A1(n2823), .A2(n2204), .ZN(n2205) );
  NOR2_X1 U2374 ( .A1(n2206), .A2(n2205), .ZN(n2207) );
  NAND2_X1 U2375 ( .A1(n2208), .A2(n2207), .ZN(n2209) );
  NOR2_X1 U2376 ( .A1(n2210), .A2(n2209), .ZN(n2211) );
  NAND2_X1 U2377 ( .A1(n2212), .A2(n2211), .ZN(N379) );
  NOR2_X1 U2378 ( .A1(n2815), .A2(n2708), .ZN(n2213) );
  NOR2_X1 U2379 ( .A1(n2214), .A2(n2213), .ZN(n2217) );
  NOR2_X1 U2380 ( .A1(n2816), .A2(SI[0]), .ZN(n2215) );
  NAND2_X1 U2381 ( .A1(n2640), .A2(n2215), .ZN(n2216) );
  NAND2_X1 U2382 ( .A1(n2217), .A2(n2216), .ZN(n2224) );
  NAND2_X1 U2383 ( .A1(SI[5]), .A2(SI[2]), .ZN(n2712) );
  NAND2_X1 U2384 ( .A1(n2712), .A2(n2769), .ZN(n2218) );
  NAND2_X1 U2385 ( .A1(n2218), .A2(n2609), .ZN(n2222) );
  NOR2_X1 U2386 ( .A1(n2298), .A2(n2672), .ZN(n2219) );
  NOR2_X1 U2387 ( .A1(n2220), .A2(n2219), .ZN(n2221) );
  NAND2_X1 U2388 ( .A1(n2222), .A2(n2221), .ZN(n2223) );
  NOR2_X1 U2389 ( .A1(n2224), .A2(n2223), .ZN(n2225) );
  NOR2_X1 U2390 ( .A1(n2828), .A2(n2225), .ZN(n2232) );
  NAND2_X1 U2391 ( .A1(n2627), .A2(n2713), .ZN(n2226) );
  NAND2_X1 U2392 ( .A1(n2504), .A2(n2226), .ZN(n2229) );
  MUX2_X1 U2393 ( .A(n2651), .B(n2227), .S(n2813), .Z(n2228) );
  NOR2_X1 U2394 ( .A1(n2229), .A2(n2228), .ZN(n2230) );
  NOR2_X1 U2395 ( .A1(n2230), .A2(n2563), .ZN(n2231) );
  NOR2_X1 U2396 ( .A1(n2232), .A2(n2231), .ZN(n2312) );
  NAND2_X1 U2397 ( .A1(n2753), .A2(n2651), .ZN(n2237) );
  NAND2_X1 U2398 ( .A1(n2417), .A2(n2813), .ZN(n2233) );
  NOR2_X1 U2399 ( .A1(n2635), .A2(n2233), .ZN(n2234) );
  NOR2_X1 U2400 ( .A1(n2235), .A2(n2234), .ZN(n2236) );
  NAND2_X1 U2401 ( .A1(n2237), .A2(n2236), .ZN(n2239) );
  NAND2_X1 U2402 ( .A1(SI[3]), .A2(n2813), .ZN(n2777) );
  NOR2_X1 U2403 ( .A1(n2777), .A2(n2631), .ZN(n2238) );
  NOR2_X1 U2404 ( .A1(n2239), .A2(n2238), .ZN(n2258) );
  NOR2_X1 U2405 ( .A1(n2707), .A2(n2713), .ZN(n2240) );
  NOR2_X1 U2406 ( .A1(n2241), .A2(n2240), .ZN(n2248) );
  NOR2_X1 U2407 ( .A1(n2709), .A2(n2242), .ZN(n2561) );
  NOR2_X1 U2408 ( .A1(SI[5]), .A2(n2442), .ZN(n2243) );
  NOR2_X1 U2409 ( .A1(n2561), .A2(n2243), .ZN(n2244) );
  NOR2_X1 U2410 ( .A1(SI[0]), .A2(n2244), .ZN(n2246) );
  NOR2_X1 U2411 ( .A1(n2615), .A2(n2442), .ZN(n2245) );
  NOR2_X1 U2412 ( .A1(n2246), .A2(n2245), .ZN(n2247) );
  NAND2_X1 U2413 ( .A1(n2248), .A2(n2247), .ZN(n2250) );
  NOR2_X1 U2414 ( .A1(n2376), .A2(n2769), .ZN(n2249) );
  NOR2_X1 U2415 ( .A1(n2250), .A2(n2249), .ZN(n2251) );
  NOR2_X1 U2416 ( .A1(n2437), .A2(n2251), .ZN(n2256) );
  MUX2_X1 U2417 ( .A(n2252), .B(n2651), .S(n2813), .Z(n2253) );
  NOR2_X1 U2418 ( .A1(n2505), .A2(n2253), .ZN(n2254) );
  NOR2_X1 U2419 ( .A1(n2254), .A2(n2785), .ZN(n2255) );
  NOR2_X1 U2420 ( .A1(n2256), .A2(n2255), .ZN(n2257) );
  NAND2_X1 U2421 ( .A1(n2258), .A2(n2257), .ZN(n2310) );
  NOR2_X1 U2422 ( .A1(n2672), .A2(n2430), .ZN(n2540) );
  NOR2_X1 U2423 ( .A1(n2261), .A2(n2640), .ZN(n2259) );
  NOR2_X1 U2424 ( .A1(n2533), .A2(n2259), .ZN(n2260) );
  NOR2_X1 U2425 ( .A1(n2540), .A2(n2260), .ZN(n2263) );
  NAND2_X1 U2426 ( .A1(n2261), .A2(n2661), .ZN(n2262) );
  NAND2_X1 U2427 ( .A1(n2263), .A2(n2262), .ZN(n2264) );
  NAND2_X1 U2428 ( .A1(n2719), .A2(n2264), .ZN(n2276) );
  NAND2_X1 U2429 ( .A1(n2417), .A2(n2789), .ZN(n2273) );
  NAND2_X1 U2430 ( .A1(n2661), .A2(n2720), .ZN(n2752) );
  NOR2_X1 U2431 ( .A1(n2315), .A2(n2777), .ZN(n2266) );
  NAND2_X1 U2432 ( .A1(n2772), .A2(n2796), .ZN(n2645) );
  NOR2_X1 U2433 ( .A1(n2645), .A2(n2791), .ZN(n2265) );
  NOR2_X1 U2434 ( .A1(n2266), .A2(n2265), .ZN(n2267) );
  NAND2_X1 U2435 ( .A1(n2752), .A2(n2267), .ZN(n2271) );
  NAND2_X1 U2436 ( .A1(SI[4]), .A2(n2725), .ZN(n2268) );
  NAND2_X1 U2437 ( .A1(n2462), .A2(n2268), .ZN(n2269) );
  NOR2_X1 U2438 ( .A1(n2635), .A2(n2269), .ZN(n2270) );
  NOR2_X1 U2439 ( .A1(n2271), .A2(n2270), .ZN(n2272) );
  NAND2_X1 U2440 ( .A1(n2273), .A2(n2272), .ZN(n2274) );
  NAND2_X1 U2441 ( .A1(n2274), .A2(SI[0]), .ZN(n2275) );
  NAND2_X1 U2442 ( .A1(n2276), .A2(n2275), .ZN(n2281) );
  NOR2_X1 U2443 ( .A1(n2816), .A2(n2786), .ZN(n2278) );
  NOR2_X1 U2444 ( .A1(n2725), .A2(n2817), .ZN(n2277) );
  NOR2_X1 U2445 ( .A1(n2278), .A2(n2277), .ZN(n2279) );
  NOR2_X1 U2446 ( .A1(n2815), .A2(n2279), .ZN(n2280) );
  NOR2_X1 U2447 ( .A1(n2281), .A2(n2280), .ZN(n2308) );
  NOR2_X1 U2448 ( .A1(n2791), .A2(n2713), .ZN(n2383) );
  NOR2_X1 U2449 ( .A1(n2694), .A2(n2383), .ZN(n2282) );
  NOR2_X1 U2450 ( .A1(n2779), .A2(n2282), .ZN(n2283) );
  NAND2_X1 U2451 ( .A1(SI[2]), .A2(n2283), .ZN(n2286) );
  NAND2_X1 U2452 ( .A1(n2736), .A2(n2533), .ZN(n2284) );
  NAND2_X1 U2453 ( .A1(n2773), .A2(n2284), .ZN(n2285) );
  NAND2_X1 U2454 ( .A1(n2286), .A2(n2285), .ZN(n2306) );
  NOR2_X1 U2455 ( .A1(n2778), .A2(n2570), .ZN(n2774) );
  NAND2_X1 U2456 ( .A1(n2774), .A2(n2760), .ZN(n2459) );
  NOR2_X1 U2457 ( .A1(n2442), .A2(n2459), .ZN(n2686) );
  NOR2_X1 U2458 ( .A1(n2823), .A2(n2778), .ZN(n2287) );
  NAND2_X1 U2459 ( .A1(SI[6]), .A2(n2287), .ZN(n2288) );
  NOR2_X1 U2460 ( .A1(SI[0]), .A2(n2288), .ZN(n2289) );
  NOR2_X1 U2461 ( .A1(n2686), .A2(n2289), .ZN(n2304) );
  NOR2_X1 U2462 ( .A1(SI[3]), .A2(n2761), .ZN(n2458) );
  NAND2_X1 U2463 ( .A1(n2458), .A2(n2672), .ZN(n2297) );
  NAND2_X1 U2464 ( .A1(n2317), .A2(n2290), .ZN(n2293) );
  NAND2_X1 U2465 ( .A1(n2624), .A2(n2291), .ZN(n2292) );
  NAND2_X1 U2466 ( .A1(n2293), .A2(n2292), .ZN(n2295) );
  NOR2_X1 U2467 ( .A1(n2616), .A2(n2642), .ZN(n2294) );
  NOR2_X1 U2468 ( .A1(n2295), .A2(n2294), .ZN(n2296) );
  NAND2_X1 U2469 ( .A1(n2297), .A2(n2296), .ZN(n2302) );
  NOR2_X1 U2470 ( .A1(n2519), .A2(n2707), .ZN(n2438) );
  NOR2_X1 U2471 ( .A1(n2298), .A2(n2315), .ZN(n2299) );
  NOR2_X1 U2472 ( .A1(n2438), .A2(n2299), .ZN(n2300) );
  NOR2_X1 U2473 ( .A1(n2723), .A2(n2300), .ZN(n2301) );
  NOR2_X1 U2474 ( .A1(n2302), .A2(n2301), .ZN(n2303) );
  NAND2_X1 U2475 ( .A1(n2304), .A2(n2303), .ZN(n2305) );
  NOR2_X1 U2476 ( .A1(n2306), .A2(n2305), .ZN(n2307) );
  NAND2_X1 U2477 ( .A1(n2308), .A2(n2307), .ZN(n2309) );
  NOR2_X1 U2478 ( .A1(n2310), .A2(n2309), .ZN(n2311) );
  NAND2_X1 U2479 ( .A1(n2312), .A2(n2311), .ZN(N470) );
  NAND2_X1 U2480 ( .A1(n2734), .A2(n2609), .ZN(n2323) );
  NAND2_X1 U2481 ( .A1(n2766), .A2(n2313), .ZN(n2371) );
  AND2_X1 U2482 ( .A1(n2571), .A2(n2371), .ZN(n2314) );
  NOR2_X1 U2483 ( .A1(SI[1]), .A2(n2314), .ZN(n2321) );
  NAND2_X1 U2484 ( .A1(n2315), .A2(n2519), .ZN(n2316) );
  NAND2_X1 U2485 ( .A1(n2316), .A2(n2682), .ZN(n2319) );
  NAND2_X1 U2486 ( .A1(n2624), .A2(n2317), .ZN(n2318) );
  NAND2_X1 U2487 ( .A1(n2319), .A2(n2318), .ZN(n2320) );
  NOR2_X1 U2488 ( .A1(n2321), .A2(n2320), .ZN(n2322) );
  NAND2_X1 U2489 ( .A1(n2323), .A2(n2322), .ZN(n2324) );
  NAND2_X1 U2490 ( .A1(n2324), .A2(n2772), .ZN(n2339) );
  NAND2_X1 U2491 ( .A1(n2642), .A2(n2498), .ZN(n2326) );
  NAND2_X1 U2492 ( .A1(n2708), .A2(n2672), .ZN(n2325) );
  NAND2_X1 U2493 ( .A1(n2326), .A2(n2325), .ZN(n2334) );
  NOR2_X1 U2494 ( .A1(n2708), .A2(n2707), .ZN(n2328) );
  NOR2_X1 U2495 ( .A1(n2742), .A2(n2723), .ZN(n2327) );
  NOR2_X1 U2496 ( .A1(n2328), .A2(n2327), .ZN(n2329) );
  NOR2_X1 U2497 ( .A1(n2329), .A2(n2779), .ZN(n2332) );
  NOR2_X1 U2498 ( .A1(n2677), .A2(n2330), .ZN(n2331) );
  NOR2_X1 U2499 ( .A1(n2332), .A2(n2331), .ZN(n2333) );
  NAND2_X1 U2500 ( .A1(n2334), .A2(n2333), .ZN(n2337) );
  NOR2_X1 U2501 ( .A1(n2417), .A2(n2674), .ZN(n2335) );
  NOR2_X1 U2502 ( .A1(n2577), .A2(n2335), .ZN(n2336) );
  NOR2_X1 U2503 ( .A1(n2337), .A2(n2336), .ZN(n2338) );
  NAND2_X1 U2504 ( .A1(n2339), .A2(n2338), .ZN(n2382) );
  NAND2_X1 U2505 ( .A1(n2737), .A2(n2694), .ZN(n2343) );
  NOR2_X1 U2506 ( .A1(n2709), .A2(n2376), .ZN(n2341) );
  NOR2_X1 U2507 ( .A1(n2810), .A2(n2736), .ZN(n2340) );
  NOR2_X1 U2508 ( .A1(n2341), .A2(n2340), .ZN(n2342) );
  NAND2_X1 U2509 ( .A1(n2343), .A2(n2342), .ZN(n2345) );
  NOR2_X1 U2510 ( .A1(n2563), .A2(n2672), .ZN(n2344) );
  NOR2_X1 U2511 ( .A1(n2345), .A2(n2344), .ZN(n2350) );
  AND2_X1 U2512 ( .A1(n2395), .A2(n2346), .ZN(n2348) );
  NOR2_X1 U2513 ( .A1(n2742), .A2(n2780), .ZN(n2347) );
  NOR2_X1 U2514 ( .A1(n2348), .A2(n2347), .ZN(n2349) );
  NAND2_X1 U2515 ( .A1(n2350), .A2(n2349), .ZN(n2351) );
  NAND2_X1 U2516 ( .A1(n2351), .A2(n2641), .ZN(n2380) );
  NAND2_X1 U2517 ( .A1(n2624), .A2(n2690), .ZN(n2375) );
  NAND2_X1 U2518 ( .A1(n2724), .A2(n2736), .ZN(n2352) );
  NAND2_X1 U2519 ( .A1(n2352), .A2(n2611), .ZN(n2367) );
  NAND2_X1 U2520 ( .A1(n2694), .A2(n2753), .ZN(n2363) );
  NAND2_X1 U2521 ( .A1(n2809), .A2(SI[1]), .ZN(n2353) );
  NAND2_X1 U2522 ( .A1(n2353), .A2(n2533), .ZN(n2354) );
  NAND2_X1 U2523 ( .A1(n2354), .A2(n2612), .ZN(n2358) );
  NOR2_X1 U2524 ( .A1(n2818), .A2(n2713), .ZN(n2355) );
  NAND2_X1 U2525 ( .A1(n2356), .A2(n2355), .ZN(n2357) );
  NAND2_X1 U2526 ( .A1(n2358), .A2(n2357), .ZN(n2361) );
  NOR2_X1 U2527 ( .A1(n2359), .A2(n2778), .ZN(n2360) );
  NOR2_X1 U2528 ( .A1(n2361), .A2(n2360), .ZN(n2362) );
  NAND2_X1 U2529 ( .A1(n2363), .A2(n2362), .ZN(n2365) );
  NOR2_X1 U2530 ( .A1(n2712), .A2(n2672), .ZN(n2364) );
  NOR2_X1 U2531 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  NAND2_X1 U2532 ( .A1(n2367), .A2(n2366), .ZN(n2368) );
  NAND2_X1 U2533 ( .A1(n2719), .A2(n2368), .ZN(n2370) );
  NAND2_X1 U2534 ( .A1(SI[3]), .A2(n2674), .ZN(n2369) );
  NAND2_X1 U2535 ( .A1(n2370), .A2(n2369), .ZN(n2373) );
  NOR2_X1 U2536 ( .A1(n2371), .A2(n2713), .ZN(n2372) );
  NOR2_X1 U2537 ( .A1(n2373), .A2(n2372), .ZN(n2374) );
  NAND2_X1 U2538 ( .A1(n2375), .A2(n2374), .ZN(n2378) );
  NOR2_X1 U2539 ( .A1(n2576), .A2(n2376), .ZN(n2377) );
  NOR2_X1 U2540 ( .A1(n2378), .A2(n2377), .ZN(n2379) );
  NAND2_X1 U2541 ( .A1(n2380), .A2(n2379), .ZN(n2381) );
  NOR2_X1 U2542 ( .A1(n2382), .A2(n2381), .ZN(n2427) );
  NOR2_X1 U2543 ( .A1(SI[4]), .A2(n2401), .ZN(n2415) );
  NAND2_X1 U2544 ( .A1(n2609), .A2(n2415), .ZN(n2467) );
  NAND2_X1 U2545 ( .A1(n2766), .A2(n2383), .ZN(n2385) );
  NAND2_X1 U2546 ( .A1(n2651), .A2(n2630), .ZN(n2384) );
  NAND2_X1 U2547 ( .A1(n2385), .A2(n2384), .ZN(n2387) );
  NOR2_X1 U2548 ( .A1(n2723), .A2(n2429), .ZN(n2386) );
  NOR2_X1 U2549 ( .A1(n2387), .A2(n2386), .ZN(n2388) );
  NAND2_X1 U2550 ( .A1(n2467), .A2(n2388), .ZN(n2389) );
  NAND2_X1 U2551 ( .A1(n2389), .A2(SI[2]), .ZN(n2399) );
  NAND2_X1 U2552 ( .A1(n2688), .A2(n2647), .ZN(n2394) );
  NAND2_X1 U2553 ( .A1(n2651), .A2(n2609), .ZN(n2391) );
  NAND2_X1 U2554 ( .A1(n2505), .A2(n2630), .ZN(n2390) );
  NAND2_X1 U2555 ( .A1(n2391), .A2(n2390), .ZN(n2392) );
  NAND2_X1 U2556 ( .A1(n2760), .A2(n2392), .ZN(n2393) );
  NAND2_X1 U2557 ( .A1(n2394), .A2(n2393), .ZN(n2397) );
  NAND2_X1 U2558 ( .A1(n2395), .A2(n2750), .ZN(n2700) );
  NOR2_X1 U2559 ( .A1(n2616), .A2(n2700), .ZN(n2396) );
  NOR2_X1 U2560 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  NAND2_X1 U2561 ( .A1(n2399), .A2(n2398), .ZN(n2425) );
  NAND2_X1 U2562 ( .A1(n2767), .A2(n2438), .ZN(n2406) );
  NOR2_X1 U2563 ( .A1(SI[3]), .A2(n2400), .ZN(n2594) );
  NOR2_X1 U2564 ( .A1(n2401), .A2(n2630), .ZN(n2402) );
  NOR2_X1 U2565 ( .A1(n2594), .A2(n2402), .ZN(n2403) );
  NOR2_X1 U2566 ( .A1(n2403), .A2(SI[6]), .ZN(n2404) );
  NAND2_X1 U2567 ( .A1(n2789), .A2(n2404), .ZN(n2405) );
  NAND2_X1 U2568 ( .A1(n2406), .A2(n2405), .ZN(n2411) );
  NOR2_X1 U2569 ( .A1(n2407), .A2(n2742), .ZN(n2408) );
  NOR2_X1 U2570 ( .A1(n2535), .A2(n2408), .ZN(n2409) );
  NOR2_X1 U2571 ( .A1(n2409), .A2(n2725), .ZN(n2410) );
  NOR2_X1 U2572 ( .A1(n2411), .A2(n2410), .ZN(n2423) );
  NOR2_X1 U2573 ( .A1(n2412), .A2(n2777), .ZN(n2574) );
  NOR2_X1 U2574 ( .A1(n2498), .A2(n2563), .ZN(n2413) );
  NOR2_X1 U2575 ( .A1(n2574), .A2(n2413), .ZN(n2414) );
  NOR2_X1 U2576 ( .A1(n2630), .A2(n2414), .ZN(n2421) );
  NAND2_X1 U2577 ( .A1(n2415), .A2(n2630), .ZN(n2416) );
  NAND2_X1 U2578 ( .A1(n2625), .A2(n2416), .ZN(n2418) );
  NOR2_X1 U2579 ( .A1(n2418), .A2(n2417), .ZN(n2419) );
  NOR2_X1 U2580 ( .A1(n2635), .A2(n2419), .ZN(n2420) );
  NOR2_X1 U2581 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  NAND2_X1 U2582 ( .A1(n2423), .A2(n2422), .ZN(n2424) );
  NOR2_X1 U2583 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  NAND2_X1 U2584 ( .A1(n2427), .A2(n2426), .ZN(N563) );
  NAND2_X1 U2585 ( .A1(n2712), .A2(n2823), .ZN(n2428) );
  NAND2_X1 U2586 ( .A1(n2428), .A2(n2641), .ZN(n2433) );
  NOR2_X1 U2587 ( .A1(SI[3]), .A2(n2429), .ZN(n2689) );
  NOR2_X1 U2588 ( .A1(n2430), .A2(n2570), .ZN(n2431) );
  NOR2_X1 U2589 ( .A1(n2689), .A2(n2431), .ZN(n2432) );
  NAND2_X1 U2590 ( .A1(n2433), .A2(n2432), .ZN(n2436) );
  NOR2_X1 U2591 ( .A1(n2647), .A2(n2492), .ZN(n2434) );
  NOR2_X1 U2592 ( .A1(SI[2]), .A2(n2434), .ZN(n2435) );
  NOR2_X1 U2593 ( .A1(n2436), .A2(n2435), .ZN(n2440) );
  NOR2_X1 U2594 ( .A1(n2437), .A2(n2615), .ZN(n2483) );
  NOR2_X1 U2595 ( .A1(n2438), .A2(n2483), .ZN(n2439) );
  NAND2_X1 U2596 ( .A1(n2440), .A2(n2439), .ZN(n2441) );
  NAND2_X1 U2597 ( .A1(n2688), .A2(n2441), .ZN(n2451) );
  NAND2_X1 U2598 ( .A1(n2766), .A2(n2540), .ZN(n2445) );
  NAND2_X1 U2599 ( .A1(n2442), .A2(n2713), .ZN(n2443) );
  NAND2_X1 U2600 ( .A1(n2690), .A2(n2443), .ZN(n2444) );
  NAND2_X1 U2601 ( .A1(n2445), .A2(n2444), .ZN(n2449) );
  NAND2_X1 U2602 ( .A1(n2790), .A2(n2446), .ZN(n2447) );
  NOR2_X1 U2603 ( .A1(SI[1]), .A2(n2447), .ZN(n2448) );
  NOR2_X1 U2604 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  NAND2_X1 U2605 ( .A1(n2451), .A2(n2450), .ZN(n2457) );
  NAND2_X1 U2606 ( .A1(n2766), .A2(n2609), .ZN(n2693) );
  NAND2_X1 U2607 ( .A1(n2761), .A2(n2693), .ZN(n2454) );
  NOR2_X1 U2608 ( .A1(n2452), .A2(n2813), .ZN(n2453) );
  NOR2_X1 U2609 ( .A1(n2454), .A2(n2453), .ZN(n2455) );
  NOR2_X1 U2610 ( .A1(n2823), .A2(n2455), .ZN(n2456) );
  NOR2_X1 U2611 ( .A1(n2457), .A2(n2456), .ZN(n2530) );
  NOR2_X1 U2612 ( .A1(n2687), .A2(n2458), .ZN(n2460) );
  NAND2_X1 U2613 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  NAND2_X1 U2614 ( .A1(SI[0]), .A2(n2461), .ZN(n2516) );
  NOR2_X1 U2615 ( .A1(SI[3]), .A2(n2462), .ZN(n2463) );
  NOR2_X1 U2616 ( .A1(n2790), .A2(n2463), .ZN(n2464) );
  NOR2_X1 U2617 ( .A1(n2791), .A2(n2464), .ZN(n2465) );
  NAND2_X1 U2618 ( .A1(n2624), .A2(n2465), .ZN(n2466) );
  NAND2_X1 U2619 ( .A1(n2467), .A2(n2466), .ZN(n2469) );
  NOR2_X1 U2620 ( .A1(n2725), .A2(n2742), .ZN(n2468) );
  MUX2_X1 U2621 ( .A(n2469), .B(n2468), .S(SI[2]), .Z(n2471) );
  NOR2_X1 U2622 ( .A1(n2813), .A2(n2576), .ZN(n2470) );
  NOR2_X1 U2623 ( .A1(n2471), .A2(n2470), .ZN(n2479) );
  NOR2_X1 U2624 ( .A1(n2778), .A2(SI[1]), .ZN(n2473) );
  NOR2_X1 U2625 ( .A1(n2815), .A2(n2780), .ZN(n2472) );
  NOR2_X1 U2626 ( .A1(n2473), .A2(n2472), .ZN(n2476) );
  NOR2_X1 U2627 ( .A1(n2810), .A2(SI[0]), .ZN(n2474) );
  NAND2_X1 U2628 ( .A1(n2661), .A2(n2474), .ZN(n2475) );
  NAND2_X1 U2629 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  NAND2_X1 U2630 ( .A1(n2719), .A2(n2477), .ZN(n2478) );
  NAND2_X1 U2631 ( .A1(n2479), .A2(n2478), .ZN(n2514) );
  NOR2_X1 U2632 ( .A1(n2810), .A2(n2828), .ZN(n2480) );
  NOR2_X1 U2633 ( .A1(n2719), .A2(n2480), .ZN(n2481) );
  NOR2_X1 U2634 ( .A1(n2769), .A2(n2481), .ZN(n2482) );
  NOR2_X1 U2635 ( .A1(n2483), .A2(n2482), .ZN(n2484) );
  NAND2_X1 U2636 ( .A1(n2761), .A2(n2484), .ZN(n2485) );
  NAND2_X1 U2637 ( .A1(n2485), .A2(n2767), .ZN(n2512) );
  NOR2_X1 U2638 ( .A1(n2577), .A2(n2615), .ZN(n2487) );
  NOR2_X1 U2639 ( .A1(n2707), .A2(n2817), .ZN(n2486) );
  NOR2_X1 U2640 ( .A1(n2487), .A2(n2486), .ZN(n2490) );
  NOR2_X1 U2641 ( .A1(n2616), .A2(n2824), .ZN(n2488) );
  NAND2_X1 U2642 ( .A1(n2661), .A2(n2488), .ZN(n2489) );
  NAND2_X1 U2643 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U2644 ( .A1(n2641), .A2(n2491), .ZN(n2502) );
  NAND2_X1 U2645 ( .A1(n2493), .A2(n2492), .ZN(n2497) );
  NOR2_X1 U2646 ( .A1(n2577), .A2(n2700), .ZN(n2495) );
  NOR2_X1 U2647 ( .A1(n2780), .A2(n2625), .ZN(n2494) );
  NOR2_X1 U2648 ( .A1(n2495), .A2(n2494), .ZN(n2496) );
  NAND2_X1 U2649 ( .A1(n2497), .A2(n2496), .ZN(n2500) );
  NOR2_X1 U2650 ( .A1(n2498), .A2(SI[0]), .ZN(n2499) );
  NOR2_X1 U2651 ( .A1(n2500), .A2(n2499), .ZN(n2501) );
  NAND2_X1 U2652 ( .A1(n2502), .A2(n2501), .ZN(n2510) );
  NAND2_X1 U2653 ( .A1(SI[0]), .A2(n2674), .ZN(n2503) );
  NAND2_X1 U2654 ( .A1(n2504), .A2(n2503), .ZN(n2507) );
  MUX2_X1 U2655 ( .A(n2505), .B(n2651), .S(n2813), .Z(n2506) );
  NOR2_X1 U2656 ( .A1(n2507), .A2(n2506), .ZN(n2508) );
  NOR2_X1 U2657 ( .A1(n2635), .A2(n2508), .ZN(n2509) );
  NOR2_X1 U2658 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  NAND2_X1 U2659 ( .A1(n2512), .A2(n2511), .ZN(n2513) );
  NOR2_X1 U2660 ( .A1(n2514), .A2(n2513), .ZN(n2515) );
  NAND2_X1 U2661 ( .A1(n2516), .A2(n2515), .ZN(n2528) );
  NAND2_X1 U2662 ( .A1(n2662), .A2(SI[1]), .ZN(n2518) );
  NAND2_X1 U2663 ( .A1(n2720), .A2(n2630), .ZN(n2517) );
  NAND2_X1 U2664 ( .A1(n2518), .A2(n2517), .ZN(n2525) );
  NAND2_X1 U2665 ( .A1(n2786), .A2(n2519), .ZN(n2520) );
  NAND2_X1 U2666 ( .A1(n2520), .A2(n2609), .ZN(n2523) );
  NOR2_X1 U2667 ( .A1(n2713), .A2(n2587), .ZN(n2521) );
  NOR2_X1 U2668 ( .A1(n2774), .A2(n2521), .ZN(n2522) );
  NAND2_X1 U2669 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  NOR2_X1 U2670 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  NOR2_X1 U2671 ( .A1(n2785), .A2(n2526), .ZN(n2527) );
  NOR2_X1 U2672 ( .A1(n2528), .A2(n2527), .ZN(n2529) );
  NAND2_X1 U2673 ( .A1(n2530), .A2(n2529), .ZN(N639) );
  NAND2_X1 U2674 ( .A1(n2737), .A2(n2595), .ZN(n2531) );
  NOR2_X1 U2675 ( .A1(SI[1]), .A2(n2531), .ZN(n2532) );
  NAND2_X1 U2676 ( .A1(n2532), .A2(SI[7]), .ZN(n2537) );
  NOR2_X1 U2677 ( .A1(n2769), .A2(n2533), .ZN(n2534) );
  NOR2_X1 U2678 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  NAND2_X1 U2679 ( .A1(n2537), .A2(n2536), .ZN(n2539) );
  NAND2_X1 U2680 ( .A1(n2539), .A2(n2538), .ZN(n2550) );
  NAND2_X1 U2681 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  NAND2_X1 U2682 ( .A1(n2543), .A2(n2542), .ZN(n2548) );
  NOR2_X1 U2683 ( .A1(n2545), .A2(n2544), .ZN(n2546) );
  NOR2_X1 U2684 ( .A1(n2724), .A2(n2546), .ZN(n2547) );
  NOR2_X1 U2685 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  NAND2_X1 U2686 ( .A1(n2550), .A2(n2549), .ZN(n2552) );
  NOR2_X1 U2687 ( .A1(n2673), .A2(n2732), .ZN(n2551) );
  NOR2_X1 U2688 ( .A1(n2552), .A2(n2551), .ZN(n2671) );
  NAND2_X1 U2689 ( .A1(n2824), .A2(n2818), .ZN(n2553) );
  NAND2_X1 U2690 ( .A1(n2553), .A2(n2679), .ZN(n2558) );
  NOR2_X1 U2691 ( .A1(n2694), .A2(n2792), .ZN(n2554) );
  NAND2_X1 U2692 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  NAND2_X1 U2693 ( .A1(n2688), .A2(n2556), .ZN(n2557) );
  NAND2_X1 U2694 ( .A1(n2558), .A2(n2557), .ZN(n2568) );
  AND2_X1 U2695 ( .A1(n2559), .A2(n2643), .ZN(n2560) );
  NOR2_X1 U2696 ( .A1(n2561), .A2(n2560), .ZN(n2566) );
  NOR2_X1 U2697 ( .A1(n2699), .A2(n2562), .ZN(n2715) );
  NOR2_X1 U2698 ( .A1(n2724), .A2(n2563), .ZN(n2564) );
  NOR2_X1 U2699 ( .A1(n2715), .A2(n2564), .ZN(n2565) );
  NAND2_X1 U2700 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  NOR2_X1 U2701 ( .A1(n2568), .A2(n2567), .ZN(n2569) );
  NOR2_X1 U2702 ( .A1(n2570), .A2(n2569), .ZN(n2593) );
  NOR2_X1 U2703 ( .A1(n2572), .A2(n2571), .ZN(n2573) );
  NOR2_X1 U2704 ( .A1(n2574), .A2(n2573), .ZN(n2591) );
  NAND2_X1 U2705 ( .A1(n2767), .A2(n2754), .ZN(n2585) );
  NAND2_X1 U2706 ( .A1(n2789), .A2(n2627), .ZN(n2581) );
  NOR2_X1 U2707 ( .A1(n2575), .A2(n2817), .ZN(n2579) );
  NOR2_X1 U2708 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
  NOR2_X1 U2709 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  NAND2_X1 U2710 ( .A1(n2581), .A2(n2580), .ZN(n2583) );
  NOR2_X1 U2711 ( .A1(n2625), .A2(n2672), .ZN(n2582) );
  NOR2_X1 U2712 ( .A1(n2583), .A2(n2582), .ZN(n2584) );
  NAND2_X1 U2713 ( .A1(n2585), .A2(n2584), .ZN(n2589) );
  NAND2_X1 U2714 ( .A1(n2688), .A2(n2694), .ZN(n2586) );
  NOR2_X1 U2715 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  NOR2_X1 U2716 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  NAND2_X1 U2717 ( .A1(n2591), .A2(n2590), .ZN(n2592) );
  NOR2_X1 U2718 ( .A1(n2593), .A2(n2592), .ZN(n2639) );
  NAND2_X1 U2719 ( .A1(n2594), .A2(n2767), .ZN(n2607) );
  NAND2_X1 U2720 ( .A1(n2595), .A2(n2643), .ZN(n2597) );
  NAND2_X1 U2721 ( .A1(n2640), .A2(n2789), .ZN(n2596) );
  NAND2_X1 U2722 ( .A1(n2597), .A2(n2596), .ZN(n2605) );
  NAND2_X1 U2723 ( .A1(n2724), .A2(n2780), .ZN(n2598) );
  NAND2_X1 U2724 ( .A1(n2598), .A2(n2611), .ZN(n2603) );
  NAND2_X1 U2725 ( .A1(n2635), .A2(SI[0]), .ZN(n2599) );
  NAND2_X1 U2726 ( .A1(n2599), .A2(n2777), .ZN(n2601) );
  NAND2_X1 U2727 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  NAND2_X1 U2728 ( .A1(n2603), .A2(n2602), .ZN(n2604) );
  NOR2_X1 U2729 ( .A1(n2605), .A2(n2604), .ZN(n2606) );
  NAND2_X1 U2730 ( .A1(n2607), .A2(n2606), .ZN(n2608) );
  NAND2_X1 U2731 ( .A1(n2608), .A2(n2766), .ZN(n2623) );
  NAND2_X1 U2732 ( .A1(n2707), .A2(n2818), .ZN(n2610) );
  NAND2_X1 U2733 ( .A1(n2610), .A2(n2609), .ZN(n2620) );
  NAND2_X1 U2734 ( .A1(n2767), .A2(n2611), .ZN(n2614) );
  NAND2_X1 U2735 ( .A1(n2612), .A2(n2789), .ZN(n2613) );
  NAND2_X1 U2736 ( .A1(n2614), .A2(n2613), .ZN(n2618) );
  NOR2_X1 U2737 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  NOR2_X1 U2738 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  NAND2_X1 U2739 ( .A1(n2620), .A2(n2619), .ZN(n2621) );
  NAND2_X1 U2740 ( .A1(n2641), .A2(n2621), .ZN(n2622) );
  NAND2_X1 U2741 ( .A1(n2623), .A2(n2622), .ZN(n2637) );
  NAND2_X1 U2742 ( .A1(n2624), .A2(n2750), .ZN(n2629) );
  NOR2_X1 U2743 ( .A1(n2813), .A2(n2625), .ZN(n2626) );
  NOR2_X1 U2744 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  NAND2_X1 U2745 ( .A1(n2629), .A2(n2628), .ZN(n2633) );
  NOR2_X1 U2746 ( .A1(n2631), .A2(n2630), .ZN(n2632) );
  NOR2_X1 U2747 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  NOR2_X1 U2748 ( .A1(n2635), .A2(n2634), .ZN(n2636) );
  NOR2_X1 U2749 ( .A1(n2637), .A2(n2636), .ZN(n2638) );
  NAND2_X1 U2750 ( .A1(n2639), .A2(n2638), .ZN(n2669) );
  NAND2_X1 U2751 ( .A1(n2641), .A2(n2640), .ZN(n2784) );
  NAND2_X1 U2752 ( .A1(n2784), .A2(n2642), .ZN(n2644) );
  NAND2_X1 U2753 ( .A1(n2644), .A2(n2643), .ZN(n2649) );
  NOR2_X1 U2754 ( .A1(SI[4]), .A2(n2645), .ZN(n2646) );
  NOR2_X1 U2755 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U2756 ( .A1(n2649), .A2(n2648), .ZN(n2660) );
  NAND2_X1 U2757 ( .A1(n2785), .A2(n2777), .ZN(n2650) );
  NAND2_X1 U2758 ( .A1(n2651), .A2(n2650), .ZN(n2653) );
  NAND2_X1 U2759 ( .A1(n2653), .A2(n2652), .ZN(n2656) );
  NOR2_X1 U2760 ( .A1(n2777), .A2(n2654), .ZN(n2655) );
  NOR2_X1 U2761 ( .A1(n2656), .A2(n2655), .ZN(n2657) );
  NAND2_X1 U2762 ( .A1(n2658), .A2(n2657), .ZN(n2659) );
  NOR2_X1 U2763 ( .A1(n2660), .A2(n2659), .ZN(n2667) );
  NAND2_X1 U2764 ( .A1(n2662), .A2(n2661), .ZN(n2663) );
  NAND2_X1 U2765 ( .A1(SI[0]), .A2(n2663), .ZN(n2664) );
  NOR2_X1 U2766 ( .A1(n2665), .A2(n2664), .ZN(n2666) );
  NOR2_X1 U2767 ( .A1(n2667), .A2(n2666), .ZN(n2668) );
  NOR2_X1 U2768 ( .A1(n2669), .A2(n2668), .ZN(n2670) );
  NAND2_X1 U2769 ( .A1(n2671), .A2(n2670), .ZN(N723) );
  NAND2_X1 U2770 ( .A1(n2673), .A2(n2672), .ZN(n2675) );
  NAND2_X1 U2771 ( .A1(n2675), .A2(n2674), .ZN(n2681) );
  NAND2_X1 U2772 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  NAND2_X1 U2773 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  NAND2_X1 U2774 ( .A1(n2681), .A2(n2680), .ZN(n2706) );
  NAND2_X1 U2775 ( .A1(n2760), .A2(n2682), .ZN(n2683) );
  NOR2_X1 U2776 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  NOR2_X1 U2777 ( .A1(n2686), .A2(n2685), .ZN(n2704) );
  NAND2_X1 U2778 ( .A1(n2687), .A2(n2724), .ZN(n2698) );
  NAND2_X1 U2779 ( .A1(n2689), .A2(n2688), .ZN(n2692) );
  NAND2_X1 U2780 ( .A1(n2690), .A2(n2789), .ZN(n2691) );
  NAND2_X1 U2781 ( .A1(n2692), .A2(n2691), .ZN(n2696) );
  NOR2_X1 U2782 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  NOR2_X1 U2783 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  NAND2_X1 U2784 ( .A1(n2698), .A2(n2697), .ZN(n2702) );
  NOR2_X1 U2785 ( .A1(n2700), .A2(n2699), .ZN(n2701) );
  NOR2_X1 U2786 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U2787 ( .A1(n2704), .A2(n2703), .ZN(n2705) );
  NOR2_X1 U2788 ( .A1(n2706), .A2(n2705), .ZN(n2832) );
  NOR2_X1 U2789 ( .A1(n2723), .A2(n2707), .ZN(n2711) );
  NOR2_X1 U2790 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  NOR2_X1 U2791 ( .A1(n2711), .A2(n2710), .ZN(n2717) );
  NOR2_X1 U2792 ( .A1(n2713), .A2(n2712), .ZN(n2714) );
  NOR2_X1 U2793 ( .A1(n2715), .A2(n2714), .ZN(n2716) );
  NAND2_X1 U2794 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  NAND2_X1 U2795 ( .A1(n2719), .A2(n2718), .ZN(n2808) );
  NAND2_X1 U2796 ( .A1(n2720), .A2(n2813), .ZN(n2729) );
  NAND2_X1 U2797 ( .A1(n2790), .A2(n2721), .ZN(n2722) );
  NOR2_X1 U2798 ( .A1(n2723), .A2(n2722), .ZN(n2727) );
  NOR2_X1 U2799 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  NOR2_X1 U2800 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  NAND2_X1 U2801 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  NAND2_X1 U2802 ( .A1(n2730), .A2(n2809), .ZN(n2747) );
  NAND2_X1 U2803 ( .A1(n2732), .A2(n2731), .ZN(n2733) );
  NOR2_X1 U2804 ( .A1(n2734), .A2(n2733), .ZN(n2735) );
  NOR2_X1 U2805 ( .A1(n2736), .A2(n2735), .ZN(n2745) );
  NOR2_X1 U2806 ( .A1(n2737), .A2(n2753), .ZN(n2738) );
  NOR2_X1 U2807 ( .A1(n2739), .A2(n2738), .ZN(n2740) );
  NOR2_X1 U2808 ( .A1(n2741), .A2(n2740), .ZN(n2743) );
  NOR2_X1 U2809 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  NOR2_X1 U2810 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  NAND2_X1 U2811 ( .A1(n2747), .A2(n2746), .ZN(n2806) );
  NOR2_X1 U2812 ( .A1(n2748), .A2(n2769), .ZN(n2749) );
  NAND2_X1 U2813 ( .A1(n2750), .A2(n2749), .ZN(n2751) );
  NAND2_X1 U2814 ( .A1(n2752), .A2(n2751), .ZN(n2759) );
  NAND2_X1 U2815 ( .A1(n2754), .A2(n2753), .ZN(n2757) );
  NAND2_X1 U2816 ( .A1(n2755), .A2(n2772), .ZN(n2756) );
  NAND2_X1 U2817 ( .A1(n2757), .A2(n2756), .ZN(n2758) );
  NOR2_X1 U2818 ( .A1(n2759), .A2(n2758), .ZN(n2804) );
  NOR2_X1 U2819 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  NOR2_X1 U2820 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  NOR2_X1 U2821 ( .A1(n2765), .A2(n2764), .ZN(n2771) );
  NAND2_X1 U2822 ( .A1(n2767), .A2(n2766), .ZN(n2768) );
  NOR2_X1 U2823 ( .A1(n2769), .A2(n2768), .ZN(n2770) );
  NOR2_X1 U2824 ( .A1(n2771), .A2(n2770), .ZN(n2802) );
  NAND2_X1 U2825 ( .A1(n2773), .A2(n2772), .ZN(n2776) );
  NAND2_X1 U2826 ( .A1(n2774), .A2(SI[3]), .ZN(n2775) );
  NAND2_X1 U2827 ( .A1(n2776), .A2(n2775), .ZN(n2800) );
  NOR2_X1 U2828 ( .A1(n2778), .A2(n2777), .ZN(n2782) );
  NOR2_X1 U2829 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NOR2_X1 U2830 ( .A1(n2782), .A2(n2781), .ZN(n2783) );
  NAND2_X1 U2831 ( .A1(n2784), .A2(n2783), .ZN(n2788) );
  NOR2_X1 U2832 ( .A1(n2786), .A2(n2785), .ZN(n2787) );
  NOR2_X1 U2833 ( .A1(n2788), .A2(n2787), .ZN(n2798) );
  NAND2_X1 U2834 ( .A1(n2790), .A2(n2789), .ZN(n2794) );
  NAND2_X1 U2835 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  NAND2_X1 U2836 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  NAND2_X1 U2837 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  NAND2_X1 U2838 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  NOR2_X1 U2839 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  MUX2_X1 U2840 ( .A(n2802), .B(n2801), .S(SI[0]), .Z(n2803) );
  NAND2_X1 U2841 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  NOR2_X1 U2842 ( .A1(n2806), .A2(n2805), .ZN(n2807) );
  NAND2_X1 U2843 ( .A1(n2808), .A2(n2807), .ZN(n2830) );
  NAND2_X1 U2844 ( .A1(n2810), .A2(n2809), .ZN(n2812) );
  NAND2_X1 U2845 ( .A1(n2812), .A2(n2811), .ZN(n2814) );
  NAND2_X1 U2846 ( .A1(n2814), .A2(n2813), .ZN(n2822) );
  NOR2_X1 U2847 ( .A1(n2816), .A2(n2815), .ZN(n2820) );
  NOR2_X1 U2848 ( .A1(n2818), .A2(n2817), .ZN(n2819) );
  NOR2_X1 U2849 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  NAND2_X1 U2850 ( .A1(n2822), .A2(n2821), .ZN(n2826) );
  NOR2_X1 U2851 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  NOR2_X1 U2852 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  NOR2_X1 U2853 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  NOR2_X1 U2854 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  NAND2_X1 U2855 ( .A1(n2832), .A2(n2831), .ZN(N789) );
endmodule

