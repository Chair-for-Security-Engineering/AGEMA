/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_BDDsylvan_ClockGating_d1 (X_s0, clk, X_s1, Fresh, rst, Y_s0, Y_s1, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input rst ;
    input [409:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output Synch ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_1390 ;

    /* cells in depth 0 */
    ClockGatingController #(17) cell_546 ( .clk (clk), .rst (rst), .GatedClk (signal_1390), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_136 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_554, signal_151}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_137 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_555, signal_152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_138 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_557, signal_153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_139 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[3]), .c ({signal_558, signal_154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_140 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[4]), .c ({signal_560, signal_155}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_141 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[5]), .c ({signal_561, signal_156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_142 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_554, signal_151}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[6]), .c ({signal_562, signal_157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_143 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_555, signal_152}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[7]), .c ({signal_563, signal_158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_144 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_554, signal_151}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[8]), .c ({signal_564, signal_159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_145 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_554, signal_151}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[9]), .c ({signal_565, signal_160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_146 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_555, signal_152}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[10]), .c ({signal_566, signal_161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_147 ( .s ({X_s1[1], X_s0[1]}), .b ({signal_555, signal_152}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[11]), .c ({signal_567, signal_162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_148 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b1}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[12]), .c ({signal_568, signal_163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_149 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b1}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[13]), .c ({signal_569, signal_164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_150 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[14]), .c ({signal_570, signal_165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_151 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[15]), .c ({signal_571, signal_166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_152 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[16]), .c ({signal_572, signal_167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_153 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[17]), .c ({signal_573, signal_168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_154 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[18]), .c ({signal_574, signal_169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_155 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[19]), .c ({signal_575, signal_170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_156 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[20]), .c ({signal_576, signal_171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_157 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[21]), .c ({signal_577, signal_172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_158 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[22]), .c ({signal_578, signal_173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_159 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[23]), .c ({signal_579, signal_174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_160 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[24]), .c ({signal_580, signal_175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_161 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[25]), .c ({signal_581, signal_176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_162 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[26]), .c ({signal_582, signal_177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_163 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[27]), .c ({signal_583, signal_178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_164 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[28]), .c ({signal_584, signal_179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_165 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[29]), .c ({signal_585, signal_180}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_166 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[30]), .c ({signal_586, signal_181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_167 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[31]), .c ({signal_587, signal_182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_168 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[32]), .c ({signal_588, signal_183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_169 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[33]), .c ({signal_589, signal_184}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_170 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[34]), .c ({signal_590, signal_185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_171 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[35]), .c ({signal_591, signal_186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_172 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[36]), .c ({signal_592, signal_187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_173 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[37]), .c ({signal_593, signal_188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_174 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[38]), .c ({signal_594, signal_189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_175 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[39]), .c ({signal_595, signal_190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_176 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[40]), .c ({signal_596, signal_191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_177 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[41]), .c ({signal_597, signal_192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_178 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[42]), .c ({signal_598, signal_193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_554, signal_151}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[43]), .c ({signal_599, signal_194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[44]), .c ({signal_600, signal_195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[45]), .c ({signal_601, signal_196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[46]), .c ({signal_602, signal_197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_183 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[47]), .c ({signal_603, signal_198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[48]), .c ({signal_604, signal_199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[49]), .c ({signal_605, signal_200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[50]), .c ({signal_606, signal_201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_187 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[51]), .c ({signal_607, signal_202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_188 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[52]), .c ({signal_608, signal_203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_189 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[53]), .c ({signal_609, signal_204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_190 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[54]), .c ({signal_610, signal_205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_191 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[55]), .c ({signal_611, signal_206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_192 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[56]), .c ({signal_612, signal_207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_193 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[57]), .c ({signal_613, signal_208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_194 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[58]), .c ({signal_614, signal_209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_195 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[59]), .c ({signal_615, signal_210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_196 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[60]), .c ({signal_616, signal_211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_197 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[61]), .c ({signal_617, signal_212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_198 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[62]), .c ({signal_618, signal_213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_199 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[63]), .c ({signal_619, signal_214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_200 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[64]), .c ({signal_620, signal_215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_201 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[65]), .c ({signal_621, signal_216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_202 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_554, signal_151}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[66]), .c ({signal_622, signal_217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_203 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[67]), .c ({signal_623, signal_218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_204 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[68]), .c ({signal_624, signal_219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_205 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[69]), .c ({signal_625, signal_220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_206 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[70]), .c ({signal_626, signal_221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_207 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[71]), .c ({signal_627, signal_222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_208 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[72]), .c ({signal_628, signal_223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_209 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[73]), .c ({signal_629, signal_224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_210 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[74]), .c ({signal_630, signal_225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_211 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[75]), .c ({signal_631, signal_226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_212 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[76]), .c ({signal_632, signal_227}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_213 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[77]), .c ({signal_633, signal_228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_214 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[78]), .c ({signal_634, signal_229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_215 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[79]), .c ({signal_635, signal_230}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_216 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[80]), .c ({signal_636, signal_231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_217 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[81]), .c ({signal_637, signal_232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_218 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[82]), .c ({signal_638, signal_233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_219 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[83]), .c ({signal_639, signal_234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_220 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[84]), .c ({signal_640, signal_235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_221 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[85]), .c ({signal_641, signal_236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_222 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[86]), .c ({signal_642, signal_237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_223 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[87]), .c ({signal_643, signal_238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_224 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[88]), .c ({signal_644, signal_239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_225 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[89]), .c ({signal_645, signal_240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_226 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[90]), .c ({signal_646, signal_241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_227 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[91]), .c ({signal_647, signal_242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_228 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[92]), .c ({signal_648, signal_243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_229 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[93]), .c ({signal_649, signal_244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_230 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[94]), .c ({signal_650, signal_245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_231 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[95]), .c ({signal_651, signal_246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_232 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[96]), .c ({signal_652, signal_247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_233 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[97]), .c ({signal_653, signal_248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_234 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[98]), .c ({signal_654, signal_249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[99]), .c ({signal_655, signal_250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[100]), .c ({signal_656, signal_251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[101]), .c ({signal_657, signal_252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[102]), .c ({signal_658, signal_253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_239 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[103]), .c ({signal_659, signal_254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[104]), .c ({signal_660, signal_255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[105]), .c ({signal_661, signal_256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[106]), .c ({signal_662, signal_257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[107]), .c ({signal_663, signal_258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_244 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[108]), .c ({signal_664, signal_259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_245 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[109]), .c ({signal_665, signal_260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_246 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_554, signal_151}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[110]), .c ({signal_666, signal_261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_247 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[111]), .c ({signal_667, signal_262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_248 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[112]), .c ({signal_668, signal_263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_249 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[113]), .c ({signal_669, signal_264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_250 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[114]), .c ({signal_670, signal_265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_251 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[115]), .c ({signal_671, signal_266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_252 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[116]), .c ({signal_672, signal_267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_253 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[117]), .c ({signal_673, signal_268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_254 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[118]), .c ({signal_674, signal_269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_255 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[119]), .c ({signal_675, signal_270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_256 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[120]), .c ({signal_676, signal_271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_257 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_558, signal_154}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[121]), .c ({signal_677, signal_272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_258 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[122]), .c ({signal_678, signal_273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_259 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[123]), .c ({signal_679, signal_274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_260 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_561, signal_156}), .clk (clk), .r (Fresh[124]), .c ({signal_680, signal_275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_261 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[125]), .c ({signal_681, signal_276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_262 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[126]), .c ({signal_682, signal_277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_263 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[127]), .c ({signal_683, signal_278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_264 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[128]), .c ({signal_684, signal_279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_265 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[129]), .c ({signal_685, signal_280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_266 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[130]), .c ({signal_686, signal_281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_267 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[131]), .c ({signal_687, signal_282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_268 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[132]), .c ({signal_688, signal_283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_269 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_563, signal_158}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[133]), .c ({signal_689, signal_284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[134]), .c ({signal_690, signal_285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_569, signal_164}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[135]), .c ({signal_691, signal_286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_272 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[136]), .c ({signal_692, signal_287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[137]), .c ({signal_693, signal_288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[138]), .c ({signal_694, signal_289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[139]), .c ({signal_695, signal_290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_571, signal_166}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[140]), .c ({signal_696, signal_291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[141]), .c ({signal_697, signal_292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[142]), .c ({signal_698, signal_293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_279 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_554, signal_151}), .clk (clk), .r (Fresh[143]), .c ({signal_699, signal_294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_280 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_562, signal_157}), .clk (clk), .r (Fresh[144]), .c ({signal_700, signal_295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_281 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_567, signal_162}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[145]), .c ({signal_701, signal_296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_282 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[146]), .c ({signal_702, signal_297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_283 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_557, signal_153}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[147]), .c ({signal_703, signal_298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_284 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_561, signal_156}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[148]), .c ({signal_704, signal_299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_285 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_554, signal_151}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[149]), .c ({signal_705, signal_300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_286 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b0}), .a ({signal_566, signal_161}), .clk (clk), .r (Fresh[150]), .c ({signal_706, signal_301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_287 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_564, signal_159}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[151]), .c ({signal_707, signal_302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_288 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_557, signal_153}), .clk (clk), .r (Fresh[152]), .c ({signal_708, signal_303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_289 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[153]), .c ({signal_709, signal_304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_290 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({signal_563, signal_158}), .clk (clk), .r (Fresh[154]), .c ({signal_710, signal_305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_291 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_562, signal_157}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[155]), .c ({signal_711, signal_306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_292 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_566, signal_161}), .a ({signal_565, signal_160}), .clk (clk), .r (Fresh[156]), .c ({signal_712, signal_307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_293 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_565, signal_160}), .a ({signal_567, signal_162}), .clk (clk), .r (Fresh[157]), .c ({signal_713, signal_308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_294 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_555, signal_152}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[158]), .c ({signal_714, signal_309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_295 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_571, signal_166}), .clk (clk), .r (Fresh[159]), .c ({signal_715, signal_310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_296 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_555, signal_152}), .a ({signal_585, signal_180}), .clk (clk), .r (Fresh[160]), .c ({signal_717, signal_311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_297 ( .s ({X_s1[2], X_s0[2]}), .b ({signal_568, signal_163}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[161]), .c ({signal_718, signal_312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_298 ( .s ({X_s1[2], X_s0[2]}), .b ({1'b0, 1'b1}), .a ({signal_569, signal_164}), .clk (clk), .r (Fresh[162]), .c ({signal_719, signal_313}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_299 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_587, signal_182}), .a ({signal_586, signal_181}), .clk (clk), .r (Fresh[163]), .c ({signal_720, signal_314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_300 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_589, signal_184}), .a ({signal_588, signal_183}), .clk (clk), .r (Fresh[164]), .c ({signal_721, signal_315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_301 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_591, signal_186}), .a ({signal_590, signal_185}), .clk (clk), .r (Fresh[165]), .c ({signal_722, signal_316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_302 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_593, signal_188}), .a ({signal_592, signal_187}), .clk (clk), .r (Fresh[166]), .c ({signal_723, signal_317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_303 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_595, signal_190}), .a ({signal_594, signal_189}), .clk (clk), .r (Fresh[167]), .c ({signal_724, signal_318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_304 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_594, signal_189}), .a ({signal_596, signal_191}), .clk (clk), .r (Fresh[168]), .c ({signal_725, signal_319}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_305 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_597, signal_192}), .a ({signal_570, signal_165}), .clk (clk), .r (Fresh[169]), .c ({signal_726, signal_320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_306 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_599, signal_194}), .a ({signal_598, signal_193}), .clk (clk), .r (Fresh[170]), .c ({signal_727, signal_321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_307 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_601, signal_196}), .a ({signal_600, signal_195}), .clk (clk), .r (Fresh[171]), .c ({signal_728, signal_322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_308 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_572, signal_167}), .a ({signal_602, signal_197}), .clk (clk), .r (Fresh[172]), .c ({signal_729, signal_323}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_309 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_604, signal_199}), .a ({signal_603, signal_198}), .clk (clk), .r (Fresh[173]), .c ({signal_730, signal_324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_310 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_605, signal_200}), .a ({signal_592, signal_187}), .clk (clk), .r (Fresh[174]), .c ({signal_731, signal_325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_311 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_607, signal_202}), .a ({signal_606, signal_201}), .clk (clk), .r (Fresh[175]), .c ({signal_732, signal_326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_312 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_609, signal_204}), .a ({signal_608, signal_203}), .clk (clk), .r (Fresh[176]), .c ({signal_733, signal_327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_313 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_611, signal_206}), .a ({signal_610, signal_205}), .clk (clk), .r (Fresh[177]), .c ({signal_734, signal_328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_314 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_613, signal_208}), .a ({signal_612, signal_207}), .clk (clk), .r (Fresh[178]), .c ({signal_735, signal_329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_315 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_615, signal_210}), .a ({signal_614, signal_209}), .clk (clk), .r (Fresh[179]), .c ({signal_736, signal_330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_316 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_617, signal_212}), .a ({signal_616, signal_211}), .clk (clk), .r (Fresh[180]), .c ({signal_737, signal_331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_317 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_598, signal_193}), .a ({signal_618, signal_213}), .clk (clk), .r (Fresh[181]), .c ({signal_738, signal_332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_318 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_620, signal_215}), .a ({signal_619, signal_214}), .clk (clk), .r (Fresh[182]), .c ({signal_739, signal_333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_319 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_622, signal_217}), .a ({signal_621, signal_216}), .clk (clk), .r (Fresh[183]), .c ({signal_740, signal_334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_320 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_624, signal_219}), .a ({signal_623, signal_218}), .clk (clk), .r (Fresh[184]), .c ({signal_741, signal_335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_321 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_625, signal_220}), .a ({signal_573, signal_168}), .clk (clk), .r (Fresh[185]), .c ({signal_742, signal_336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_322 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_627, signal_222}), .a ({signal_626, signal_221}), .clk (clk), .r (Fresh[186]), .c ({signal_743, signal_337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_323 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_629, signal_224}), .a ({signal_628, signal_223}), .clk (clk), .r (Fresh[187]), .c ({signal_744, signal_338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_324 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_631, signal_226}), .a ({signal_630, signal_225}), .clk (clk), .r (Fresh[188]), .c ({signal_745, signal_339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_325 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_632, signal_227}), .a ({signal_616, signal_211}), .clk (clk), .r (Fresh[189]), .c ({signal_746, signal_340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_326 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_592, signal_187}), .a ({signal_590, signal_185}), .clk (clk), .r (Fresh[190]), .c ({signal_747, signal_341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_327 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_634, signal_229}), .a ({signal_633, signal_228}), .clk (clk), .r (Fresh[191]), .c ({signal_748, signal_342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_328 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_635, signal_230}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[192]), .c ({signal_749, signal_343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_329 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_574, signal_169}), .a ({signal_630, signal_225}), .clk (clk), .r (Fresh[193]), .c ({signal_750, signal_344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_330 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_635, signal_230}), .a ({signal_575, signal_170}), .clk (clk), .r (Fresh[194]), .c ({signal_751, signal_345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_331 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_589, signal_184}), .a ({signal_576, signal_171}), .clk (clk), .r (Fresh[195]), .c ({signal_752, signal_346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_332 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_570, signal_165}), .a ({signal_636, signal_231}), .clk (clk), .r (Fresh[196]), .c ({signal_753, signal_347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_333 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_638, signal_233}), .a ({signal_637, signal_232}), .clk (clk), .r (Fresh[197]), .c ({signal_754, signal_348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_334 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_575, signal_170}), .a ({signal_624, signal_219}), .clk (clk), .r (Fresh[198]), .c ({signal_755, signal_349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_335 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_635, signal_230}), .a ({signal_639, signal_234}), .clk (clk), .r (Fresh[199]), .c ({signal_756, signal_350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_336 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_641, signal_236}), .a ({signal_640, signal_235}), .clk (clk), .r (Fresh[200]), .c ({signal_757, signal_351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_337 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_577, signal_172}), .a ({signal_642, signal_237}), .clk (clk), .r (Fresh[201]), .c ({signal_758, signal_352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_338 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_643, signal_238}), .a ({signal_578, signal_173}), .clk (clk), .r (Fresh[202]), .c ({signal_759, signal_353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_339 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_645, signal_240}), .a ({signal_644, signal_239}), .clk (clk), .r (Fresh[203]), .c ({signal_760, signal_354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_340 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_647, signal_242}), .a ({signal_646, signal_241}), .clk (clk), .r (Fresh[204]), .c ({signal_761, signal_355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_341 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_649, signal_244}), .a ({signal_648, signal_243}), .clk (clk), .r (Fresh[205]), .c ({signal_762, signal_356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_342 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_591, signal_186}), .a ({signal_650, signal_245}), .clk (clk), .r (Fresh[206]), .c ({signal_763, signal_357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_343 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_652, signal_247}), .a ({signal_651, signal_246}), .clk (clk), .r (Fresh[207]), .c ({signal_764, signal_358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_344 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_643, signal_238}), .a ({signal_653, signal_248}), .clk (clk), .r (Fresh[208]), .c ({signal_765, signal_359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_345 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_654, signal_249}), .a ({signal_642, signal_237}), .clk (clk), .r (Fresh[209]), .c ({signal_766, signal_360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_346 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_655, signal_250}), .a ({signal_627, signal_222}), .clk (clk), .r (Fresh[210]), .c ({signal_767, signal_361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_347 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_656, signal_251}), .a ({signal_607, signal_202}), .clk (clk), .r (Fresh[211]), .c ({signal_768, signal_362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_348 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_658, signal_253}), .a ({signal_657, signal_252}), .clk (clk), .r (Fresh[212]), .c ({signal_769, signal_363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_349 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_659, signal_254}), .a ({signal_614, signal_209}), .clk (clk), .r (Fresh[213]), .c ({signal_770, signal_364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_350 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_660, signal_255}), .a ({signal_643, signal_238}), .clk (clk), .r (Fresh[214]), .c ({signal_771, signal_365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_351 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_662, signal_257}), .a ({signal_661, signal_256}), .clk (clk), .r (Fresh[215]), .c ({signal_772, signal_366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_352 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_664, signal_259}), .a ({signal_663, signal_258}), .clk (clk), .r (Fresh[216]), .c ({signal_773, signal_367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_353 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_576, signal_171}), .a ({signal_665, signal_260}), .clk (clk), .r (Fresh[217]), .c ({signal_774, signal_368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_354 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_660, signal_255}), .a ({signal_611, signal_206}), .clk (clk), .r (Fresh[218]), .c ({signal_775, signal_369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_355 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_600, signal_195}), .a ({signal_666, signal_261}), .clk (clk), .r (Fresh[219]), .c ({signal_776, signal_370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_356 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_624, signal_219}), .a ({signal_598, signal_193}), .clk (clk), .r (Fresh[220]), .c ({signal_777, signal_371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_357 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_645, signal_240}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[221]), .c ({signal_778, signal_372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_358 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_635, signal_230}), .a ({signal_667, signal_262}), .clk (clk), .r (Fresh[222]), .c ({signal_779, signal_373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_359 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_668, signal_263}), .a ({signal_594, signal_189}), .clk (clk), .r (Fresh[223]), .c ({signal_780, signal_374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_360 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_647, signal_242}), .a ({signal_669, signal_264}), .clk (clk), .r (Fresh[224]), .c ({signal_781, signal_375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_361 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_671, signal_266}), .a ({signal_670, signal_265}), .clk (clk), .r (Fresh[225]), .c ({signal_782, signal_376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_362 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_621, signal_216}), .a ({signal_672, signal_267}), .clk (clk), .r (Fresh[226]), .c ({signal_783, signal_377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_363 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_594, signal_189}), .a ({signal_673, signal_268}), .clk (clk), .r (Fresh[227]), .c ({signal_784, signal_378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_364 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_634, signal_229}), .a ({signal_579, signal_174}), .clk (clk), .r (Fresh[228]), .c ({signal_785, signal_379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_365 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_674, signal_269}), .a ({signal_638, signal_233}), .clk (clk), .r (Fresh[229]), .c ({signal_786, signal_380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_366 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_574, signal_169}), .a ({signal_624, signal_219}), .clk (clk), .r (Fresh[230]), .c ({signal_787, signal_381}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_367 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_591, signal_186}), .a ({signal_675, signal_270}), .clk (clk), .r (Fresh[231]), .c ({signal_788, signal_382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_368 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_626, signal_221}), .a ({signal_596, signal_191}), .clk (clk), .r (Fresh[232]), .c ({signal_789, signal_383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_369 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_654, signal_249}), .a ({signal_676, signal_271}), .clk (clk), .r (Fresh[233]), .c ({signal_790, signal_384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_370 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_627, signal_222}), .a ({signal_677, signal_272}), .clk (clk), .r (Fresh[234]), .c ({signal_791, signal_385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_371 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_679, signal_274}), .a ({signal_678, signal_273}), .clk (clk), .r (Fresh[235]), .c ({signal_792, signal_386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_372 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_680, signal_275}), .a ({signal_592, signal_187}), .clk (clk), .r (Fresh[236]), .c ({signal_793, signal_387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_373 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_681, signal_276}), .a ({signal_630, signal_225}), .clk (clk), .r (Fresh[237]), .c ({signal_794, signal_388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_374 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_672, signal_267}), .a ({signal_560, signal_155}), .clk (clk), .r (Fresh[238]), .c ({signal_795, signal_389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_375 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_683, signal_278}), .a ({signal_682, signal_277}), .clk (clk), .r (Fresh[239]), .c ({signal_796, signal_390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_376 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_568, signal_163}), .a ({signal_684, signal_279}), .clk (clk), .r (Fresh[240]), .c ({signal_797, signal_391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_377 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_685, signal_280}), .a ({signal_667, signal_262}), .clk (clk), .r (Fresh[241]), .c ({signal_798, signal_392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_378 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_587, signal_182}), .a ({signal_606, signal_201}), .clk (clk), .r (Fresh[242]), .c ({signal_799, signal_393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_379 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_596, signal_191}), .a ({signal_686, signal_281}), .clk (clk), .r (Fresh[243]), .c ({signal_800, signal_394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_380 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_605, signal_200}), .a ({signal_654, signal_249}), .clk (clk), .r (Fresh[244]), .c ({signal_801, signal_395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_381 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_586, signal_181}), .a ({signal_623, signal_218}), .clk (clk), .r (Fresh[245]), .c ({signal_802, signal_396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_382 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_590, signal_185}), .a ({signal_666, signal_261}), .clk (clk), .r (Fresh[246]), .c ({signal_803, signal_397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_383 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_687, signal_282}), .a ({signal_635, signal_230}), .clk (clk), .r (Fresh[247]), .c ({signal_804, signal_398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_384 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_674, signal_269}), .a ({signal_558, signal_154}), .clk (clk), .r (Fresh[248]), .c ({signal_805, signal_399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_385 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_688, signal_283}), .a ({signal_597, signal_192}), .clk (clk), .r (Fresh[249]), .c ({signal_806, signal_400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_386 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_690, signal_285}), .a ({signal_689, signal_284}), .clk (clk), .r (Fresh[250]), .c ({signal_807, signal_401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_387 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_682, signal_277}), .a ({signal_691, signal_286}), .clk (clk), .r (Fresh[251]), .c ({signal_808, signal_402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_388 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_607, signal_202}), .a ({signal_555, signal_152}), .clk (clk), .r (Fresh[252]), .c ({signal_809, signal_403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_389 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_693, signal_288}), .a ({signal_692, signal_287}), .clk (clk), .r (Fresh[253]), .c ({signal_810, signal_404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_390 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_648, signal_243}), .a ({signal_592, signal_187}), .clk (clk), .r (Fresh[254]), .c ({signal_811, signal_405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_391 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_593, signal_188}), .a ({signal_694, signal_289}), .clk (clk), .r (Fresh[255]), .c ({signal_812, signal_406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_392 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_633, signal_228}), .a ({signal_580, signal_175}), .clk (clk), .r (Fresh[256]), .c ({signal_813, signal_407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_393 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_696, signal_291}), .a ({signal_695, signal_290}), .clk (clk), .r (Fresh[257]), .c ({signal_814, signal_408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_394 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_697, signal_292}), .a ({signal_564, signal_159}), .clk (clk), .r (Fresh[258]), .c ({signal_815, signal_409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_395 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_641, signal_236}), .a ({signal_698, signal_293}), .clk (clk), .r (Fresh[259]), .c ({signal_816, signal_410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_396 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_557, signal_153}), .a ({signal_685, signal_280}), .clk (clk), .r (Fresh[260]), .c ({signal_817, signal_411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_397 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_699, signal_294}), .a ({signal_666, signal_261}), .clk (clk), .r (Fresh[261]), .c ({signal_818, signal_412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_398 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_701, signal_296}), .a ({signal_700, signal_295}), .clk (clk), .r (Fresh[262]), .c ({signal_819, signal_413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_399 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_691, signal_286}), .a ({signal_578, signal_173}), .clk (clk), .r (Fresh[263]), .c ({signal_820, signal_414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_400 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_702, signal_297}), .a ({signal_604, signal_199}), .clk (clk), .r (Fresh[264]), .c ({signal_821, signal_415}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_401 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_692, signal_287}), .a ({signal_703, signal_298}), .clk (clk), .r (Fresh[265]), .c ({signal_822, signal_416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_402 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_699, signal_294}), .a ({signal_599, signal_194}), .clk (clk), .r (Fresh[266]), .c ({signal_823, signal_417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_403 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_705, signal_300}), .a ({signal_704, signal_299}), .clk (clk), .r (Fresh[267]), .c ({signal_824, signal_418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_404 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_642, signal_237}), .a ({signal_660, signal_255}), .clk (clk), .r (Fresh[268]), .c ({signal_825, signal_419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_405 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_601, signal_196}), .a ({signal_573, signal_168}), .clk (clk), .r (Fresh[269]), .c ({signal_826, signal_420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_406 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_706, signal_301}), .a ({signal_666, signal_261}), .clk (clk), .r (Fresh[270]), .c ({signal_827, signal_421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_407 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_581, signal_176}), .a ({signal_696, signal_291}), .clk (clk), .r (Fresh[271]), .c ({signal_828, signal_422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_408 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_682, signal_277}), .a ({signal_582, signal_177}), .clk (clk), .r (Fresh[272]), .c ({signal_829, signal_423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_409 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_707, signal_302}), .a ({signal_682, signal_277}), .clk (clk), .r (Fresh[273]), .c ({signal_830, signal_424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_410 ( .s ({X_s1[3], X_s0[3]}), .b ({1'b0, 1'b1}), .a ({signal_627, signal_222}), .clk (clk), .r (Fresh[274]), .c ({signal_831, signal_425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_411 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_708, signal_303}), .a ({signal_667, signal_262}), .clk (clk), .r (Fresh[275]), .c ({signal_832, signal_426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_412 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_709, signal_304}), .a ({signal_656, signal_251}), .clk (clk), .r (Fresh[276]), .c ({signal_833, signal_427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_413 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_561, signal_156}), .a ({signal_685, signal_280}), .clk (clk), .r (Fresh[277]), .c ({signal_834, signal_428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_414 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_710, signal_305}), .a ({signal_681, signal_276}), .clk (clk), .r (Fresh[278]), .c ({signal_835, signal_429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_415 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_703, signal_298}), .a ({signal_630, signal_225}), .clk (clk), .r (Fresh[279]), .c ({signal_836, signal_430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_416 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_711, signal_306}), .a ({signal_568, signal_163}), .clk (clk), .r (Fresh[280]), .c ({signal_837, signal_431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_417 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_583, signal_178}), .a ({signal_712, signal_307}), .clk (clk), .r (Fresh[281]), .c ({signal_838, signal_432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_418 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_713, signal_308}), .a ({signal_584, signal_179}), .clk (clk), .r (Fresh[282]), .c ({signal_839, signal_433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_419 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_714, signal_309}), .a ({signal_709, signal_304}), .clk (clk), .r (Fresh[283]), .c ({signal_840, signal_434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_420 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_715, signal_310}), .a ({signal_682, signal_277}), .clk (clk), .r (Fresh[284]), .c ({signal_841, signal_435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_421 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_621, signal_216}), .a ({signal_626, signal_221}), .clk (clk), .r (Fresh[285]), .c ({signal_842, signal_436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_422 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_701, signal_296}), .a ({signal_576, signal_171}), .clk (clk), .r (Fresh[286]), .c ({signal_843, signal_437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_423 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_718, signal_312}), .a ({signal_624, signal_219}), .clk (clk), .r (Fresh[287]), .c ({signal_844, signal_438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_424 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_616, signal_211}), .a ({signal_719, signal_313}), .clk (clk), .r (Fresh[288]), .c ({signal_845, signal_439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_425 ( .s ({X_s1[3], X_s0[3]}), .b ({signal_668, signal_263}), .a ({signal_615, signal_210}), .clk (clk), .r (Fresh[289]), .c ({signal_846, signal_440}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_426 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_721, signal_315}), .a ({signal_720, signal_314}), .clk (clk), .r (Fresh[290]), .c ({signal_848, signal_441}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_427 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_723, signal_317}), .a ({signal_722, signal_316}), .clk (clk), .r (Fresh[291]), .c ({signal_849, signal_442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_428 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_725, signal_319}), .a ({signal_724, signal_318}), .clk (clk), .r (Fresh[292]), .c ({signal_850, signal_443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_429 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_727, signal_321}), .a ({signal_726, signal_320}), .clk (clk), .r (Fresh[293]), .c ({signal_851, signal_444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_430 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_729, signal_323}), .a ({signal_728, signal_322}), .clk (clk), .r (Fresh[294]), .c ({signal_852, signal_445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_431 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_731, signal_325}), .a ({signal_730, signal_324}), .clk (clk), .r (Fresh[295]), .c ({signal_853, signal_446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_432 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_733, signal_327}), .a ({signal_732, signal_326}), .clk (clk), .r (Fresh[296]), .c ({signal_854, signal_447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_433 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_735, signal_329}), .a ({signal_734, signal_328}), .clk (clk), .r (Fresh[297]), .c ({signal_855, signal_448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_434 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_737, signal_331}), .a ({signal_736, signal_330}), .clk (clk), .r (Fresh[298]), .c ({signal_856, signal_449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_435 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_739, signal_333}), .a ({signal_738, signal_332}), .clk (clk), .r (Fresh[299]), .c ({signal_857, signal_450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_436 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_741, signal_335}), .a ({signal_740, signal_334}), .clk (clk), .r (Fresh[300]), .c ({signal_858, signal_451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_437 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_743, signal_337}), .a ({signal_742, signal_336}), .clk (clk), .r (Fresh[301]), .c ({signal_859, signal_452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_438 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_745, signal_339}), .a ({signal_744, signal_338}), .clk (clk), .r (Fresh[302]), .c ({signal_860, signal_453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_439 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_747, signal_341}), .a ({signal_746, signal_340}), .clk (clk), .r (Fresh[303]), .c ({signal_861, signal_454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_440 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_749, signal_343}), .a ({signal_748, signal_342}), .clk (clk), .r (Fresh[304]), .c ({signal_862, signal_455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_441 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_751, signal_345}), .a ({signal_750, signal_344}), .clk (clk), .r (Fresh[305]), .c ({signal_863, signal_456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_442 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_753, signal_347}), .a ({signal_752, signal_346}), .clk (clk), .r (Fresh[306]), .c ({signal_864, signal_457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_443 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_755, signal_349}), .a ({signal_754, signal_348}), .clk (clk), .r (Fresh[307]), .c ({signal_865, signal_458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_444 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_757, signal_351}), .a ({signal_756, signal_350}), .clk (clk), .r (Fresh[308]), .c ({signal_866, signal_459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_445 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_759, signal_353}), .a ({signal_758, signal_352}), .clk (clk), .r (Fresh[309]), .c ({signal_867, signal_460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_446 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_761, signal_355}), .a ({signal_760, signal_354}), .clk (clk), .r (Fresh[310]), .c ({signal_868, signal_461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_447 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_763, signal_357}), .a ({signal_762, signal_356}), .clk (clk), .r (Fresh[311]), .c ({signal_869, signal_462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_448 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_765, signal_359}), .a ({signal_764, signal_358}), .clk (clk), .r (Fresh[312]), .c ({signal_870, signal_463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_449 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_767, signal_361}), .a ({signal_766, signal_360}), .clk (clk), .r (Fresh[313]), .c ({signal_871, signal_464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_450 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_769, signal_363}), .a ({signal_768, signal_362}), .clk (clk), .r (Fresh[314]), .c ({signal_872, signal_465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_451 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_771, signal_365}), .a ({signal_770, signal_364}), .clk (clk), .r (Fresh[315]), .c ({signal_873, signal_466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_452 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_773, signal_367}), .a ({signal_772, signal_366}), .clk (clk), .r (Fresh[316]), .c ({signal_874, signal_467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_453 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_775, signal_369}), .a ({signal_774, signal_368}), .clk (clk), .r (Fresh[317]), .c ({signal_875, signal_468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_454 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_777, signal_371}), .a ({signal_776, signal_370}), .clk (clk), .r (Fresh[318]), .c ({signal_876, signal_469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_455 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_779, signal_373}), .a ({signal_778, signal_372}), .clk (clk), .r (Fresh[319]), .c ({signal_877, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_456 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_781, signal_375}), .a ({signal_780, signal_374}), .clk (clk), .r (Fresh[320]), .c ({signal_878, signal_471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_457 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_783, signal_377}), .a ({signal_782, signal_376}), .clk (clk), .r (Fresh[321]), .c ({signal_879, signal_472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_458 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_785, signal_379}), .a ({signal_784, signal_378}), .clk (clk), .r (Fresh[322]), .c ({signal_880, signal_473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_459 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_787, signal_381}), .a ({signal_786, signal_380}), .clk (clk), .r (Fresh[323]), .c ({signal_881, signal_474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_460 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_789, signal_383}), .a ({signal_788, signal_382}), .clk (clk), .r (Fresh[324]), .c ({signal_882, signal_475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_461 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_791, signal_385}), .a ({signal_790, signal_384}), .clk (clk), .r (Fresh[325]), .c ({signal_883, signal_476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_462 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_793, signal_387}), .a ({signal_792, signal_386}), .clk (clk), .r (Fresh[326]), .c ({signal_884, signal_477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_463 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_795, signal_389}), .a ({signal_794, signal_388}), .clk (clk), .r (Fresh[327]), .c ({signal_885, signal_478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_464 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_797, signal_391}), .a ({signal_796, signal_390}), .clk (clk), .r (Fresh[328]), .c ({signal_886, signal_479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_465 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_799, signal_393}), .a ({signal_798, signal_392}), .clk (clk), .r (Fresh[329]), .c ({signal_887, signal_480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_466 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_801, signal_395}), .a ({signal_800, signal_394}), .clk (clk), .r (Fresh[330]), .c ({signal_888, signal_481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_467 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_803, signal_397}), .a ({signal_802, signal_396}), .clk (clk), .r (Fresh[331]), .c ({signal_889, signal_482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_468 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_805, signal_399}), .a ({signal_804, signal_398}), .clk (clk), .r (Fresh[332]), .c ({signal_890, signal_483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_469 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_807, signal_401}), .a ({signal_806, signal_400}), .clk (clk), .r (Fresh[333]), .c ({signal_891, signal_484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_470 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_809, signal_403}), .a ({signal_808, signal_402}), .clk (clk), .r (Fresh[334]), .c ({signal_892, signal_485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_471 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_811, signal_405}), .a ({signal_810, signal_404}), .clk (clk), .r (Fresh[335]), .c ({signal_893, signal_486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_472 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_813, signal_407}), .a ({signal_812, signal_406}), .clk (clk), .r (Fresh[336]), .c ({signal_894, signal_487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_473 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_815, signal_409}), .a ({signal_814, signal_408}), .clk (clk), .r (Fresh[337]), .c ({signal_895, signal_488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_474 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_817, signal_411}), .a ({signal_816, signal_410}), .clk (clk), .r (Fresh[338]), .c ({signal_896, signal_489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_475 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_819, signal_413}), .a ({signal_818, signal_412}), .clk (clk), .r (Fresh[339]), .c ({signal_897, signal_490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_476 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_821, signal_415}), .a ({signal_820, signal_414}), .clk (clk), .r (Fresh[340]), .c ({signal_898, signal_491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_477 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_823, signal_417}), .a ({signal_822, signal_416}), .clk (clk), .r (Fresh[341]), .c ({signal_899, signal_492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_478 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_825, signal_419}), .a ({signal_824, signal_418}), .clk (clk), .r (Fresh[342]), .c ({signal_900, signal_493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_479 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_827, signal_421}), .a ({signal_826, signal_420}), .clk (clk), .r (Fresh[343]), .c ({signal_901, signal_494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_480 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_829, signal_423}), .a ({signal_828, signal_422}), .clk (clk), .r (Fresh[344]), .c ({signal_902, signal_495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_481 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_831, signal_425}), .a ({signal_830, signal_424}), .clk (clk), .r (Fresh[345]), .c ({signal_903, signal_496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_482 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_833, signal_427}), .a ({signal_832, signal_426}), .clk (clk), .r (Fresh[346]), .c ({signal_904, signal_497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_483 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_835, signal_429}), .a ({signal_834, signal_428}), .clk (clk), .r (Fresh[347]), .c ({signal_905, signal_498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_484 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_837, signal_431}), .a ({signal_836, signal_430}), .clk (clk), .r (Fresh[348]), .c ({signal_906, signal_499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_485 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_839, signal_433}), .a ({signal_838, signal_432}), .clk (clk), .r (Fresh[349]), .c ({signal_907, signal_500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_486 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_841, signal_435}), .a ({signal_840, signal_434}), .clk (clk), .r (Fresh[350]), .c ({signal_908, signal_501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_487 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_843, signal_437}), .a ({signal_842, signal_436}), .clk (clk), .r (Fresh[351]), .c ({signal_909, signal_502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_488 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_844, signal_438}), .a ({signal_717, signal_311}), .clk (clk), .r (Fresh[352]), .c ({signal_910, signal_503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_489 ( .s ({X_s1[4], X_s0[4]}), .b ({signal_846, signal_440}), .a ({signal_845, signal_439}), .clk (clk), .r (Fresh[353]), .c ({signal_911, signal_504}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_490 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_849, signal_442}), .a ({signal_848, signal_441}), .clk (clk), .r (Fresh[354]), .c ({signal_913, signal_505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_491 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_851, signal_444}), .a ({signal_850, signal_443}), .clk (clk), .r (Fresh[355]), .c ({signal_914, signal_506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_492 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_853, signal_446}), .a ({signal_852, signal_445}), .clk (clk), .r (Fresh[356]), .c ({signal_915, signal_507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_493 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_855, signal_448}), .a ({signal_854, signal_447}), .clk (clk), .r (Fresh[357]), .c ({signal_916, signal_508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_494 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_857, signal_450}), .a ({signal_856, signal_449}), .clk (clk), .r (Fresh[358]), .c ({signal_917, signal_509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_495 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_859, signal_452}), .a ({signal_858, signal_451}), .clk (clk), .r (Fresh[359]), .c ({signal_918, signal_510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_496 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_861, signal_454}), .a ({signal_860, signal_453}), .clk (clk), .r (Fresh[360]), .c ({signal_919, signal_511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_497 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_863, signal_456}), .a ({signal_862, signal_455}), .clk (clk), .r (Fresh[361]), .c ({signal_920, signal_512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_498 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_865, signal_458}), .a ({signal_864, signal_457}), .clk (clk), .r (Fresh[362]), .c ({signal_921, signal_513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_499 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_867, signal_460}), .a ({signal_866, signal_459}), .clk (clk), .r (Fresh[363]), .c ({signal_922, signal_514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_500 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_869, signal_462}), .a ({signal_868, signal_461}), .clk (clk), .r (Fresh[364]), .c ({signal_923, signal_515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_501 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_871, signal_464}), .a ({signal_870, signal_463}), .clk (clk), .r (Fresh[365]), .c ({signal_924, signal_516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_502 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_873, signal_466}), .a ({signal_872, signal_465}), .clk (clk), .r (Fresh[366]), .c ({signal_925, signal_517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_503 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_875, signal_468}), .a ({signal_874, signal_467}), .clk (clk), .r (Fresh[367]), .c ({signal_926, signal_518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_504 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_877, signal_470}), .a ({signal_876, signal_469}), .clk (clk), .r (Fresh[368]), .c ({signal_927, signal_519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_505 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_879, signal_472}), .a ({signal_878, signal_471}), .clk (clk), .r (Fresh[369]), .c ({signal_928, signal_520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_506 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_881, signal_474}), .a ({signal_880, signal_473}), .clk (clk), .r (Fresh[370]), .c ({signal_929, signal_521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_507 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_883, signal_476}), .a ({signal_882, signal_475}), .clk (clk), .r (Fresh[371]), .c ({signal_930, signal_522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_508 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_885, signal_478}), .a ({signal_884, signal_477}), .clk (clk), .r (Fresh[372]), .c ({signal_931, signal_523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_509 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_887, signal_480}), .a ({signal_886, signal_479}), .clk (clk), .r (Fresh[373]), .c ({signal_932, signal_524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_510 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_889, signal_482}), .a ({signal_888, signal_481}), .clk (clk), .r (Fresh[374]), .c ({signal_933, signal_525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_511 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_891, signal_484}), .a ({signal_890, signal_483}), .clk (clk), .r (Fresh[375]), .c ({signal_934, signal_526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_512 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_893, signal_486}), .a ({signal_892, signal_485}), .clk (clk), .r (Fresh[376]), .c ({signal_935, signal_527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_513 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_895, signal_488}), .a ({signal_894, signal_487}), .clk (clk), .r (Fresh[377]), .c ({signal_936, signal_528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_514 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_897, signal_490}), .a ({signal_896, signal_489}), .clk (clk), .r (Fresh[378]), .c ({signal_937, signal_529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_515 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_899, signal_492}), .a ({signal_898, signal_491}), .clk (clk), .r (Fresh[379]), .c ({signal_938, signal_530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_516 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_901, signal_494}), .a ({signal_900, signal_493}), .clk (clk), .r (Fresh[380]), .c ({signal_939, signal_531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_517 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_903, signal_496}), .a ({signal_902, signal_495}), .clk (clk), .r (Fresh[381]), .c ({signal_940, signal_532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_518 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_905, signal_498}), .a ({signal_904, signal_497}), .clk (clk), .r (Fresh[382]), .c ({signal_941, signal_533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_519 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_907, signal_500}), .a ({signal_906, signal_499}), .clk (clk), .r (Fresh[383]), .c ({signal_942, signal_534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_520 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_909, signal_502}), .a ({signal_908, signal_501}), .clk (clk), .r (Fresh[384]), .c ({signal_943, signal_535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_521 ( .s ({X_s1[5], X_s0[5]}), .b ({signal_911, signal_504}), .a ({signal_910, signal_503}), .clk (clk), .r (Fresh[385]), .c ({signal_944, signal_536}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_522 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_914, signal_506}), .a ({signal_913, signal_505}), .clk (clk), .r (Fresh[386]), .c ({signal_946, signal_537}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_523 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_916, signal_508}), .a ({signal_915, signal_507}), .clk (clk), .r (Fresh[387]), .c ({signal_947, signal_538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_524 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_918, signal_510}), .a ({signal_917, signal_509}), .clk (clk), .r (Fresh[388]), .c ({signal_948, signal_539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_525 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_920, signal_512}), .a ({signal_919, signal_511}), .clk (clk), .r (Fresh[389]), .c ({signal_949, signal_540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_526 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_922, signal_514}), .a ({signal_921, signal_513}), .clk (clk), .r (Fresh[390]), .c ({signal_950, signal_541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_527 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_924, signal_516}), .a ({signal_923, signal_515}), .clk (clk), .r (Fresh[391]), .c ({signal_951, signal_542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_528 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_926, signal_518}), .a ({signal_925, signal_517}), .clk (clk), .r (Fresh[392]), .c ({signal_952, signal_543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_529 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_928, signal_520}), .a ({signal_927, signal_519}), .clk (clk), .r (Fresh[393]), .c ({signal_953, signal_544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_530 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_930, signal_522}), .a ({signal_929, signal_521}), .clk (clk), .r (Fresh[394]), .c ({signal_954, signal_545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_531 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_932, signal_524}), .a ({signal_931, signal_523}), .clk (clk), .r (Fresh[395]), .c ({signal_955, signal_546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_532 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_934, signal_526}), .a ({signal_933, signal_525}), .clk (clk), .r (Fresh[396]), .c ({signal_956, signal_547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_533 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_936, signal_528}), .a ({signal_935, signal_527}), .clk (clk), .r (Fresh[397]), .c ({signal_957, signal_548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_534 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_938, signal_530}), .a ({signal_937, signal_529}), .clk (clk), .r (Fresh[398]), .c ({signal_958, signal_549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_535 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_940, signal_532}), .a ({signal_939, signal_531}), .clk (clk), .r (Fresh[399]), .c ({signal_959, signal_550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_536 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_942, signal_534}), .a ({signal_941, signal_533}), .clk (clk), .r (Fresh[400]), .c ({signal_960, signal_551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_537 ( .s ({X_s1[6], X_s0[6]}), .b ({signal_944, signal_536}), .a ({signal_943, signal_535}), .clk (clk), .r (Fresh[401]), .c ({signal_961, signal_552}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_538 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_947, signal_538}), .a ({signal_946, signal_537}), .clk (clk), .r (Fresh[402]), .c ({signal_963, signal_150}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_539 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_949, signal_540}), .a ({signal_948, signal_539}), .clk (clk), .r (Fresh[403]), .c ({signal_964, signal_149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_540 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_951, signal_542}), .a ({signal_950, signal_541}), .clk (clk), .r (Fresh[404]), .c ({signal_965, signal_148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_541 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_953, signal_544}), .a ({signal_952, signal_543}), .clk (clk), .r (Fresh[405]), .c ({signal_966, signal_147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_542 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_955, signal_546}), .a ({signal_954, signal_545}), .clk (clk), .r (Fresh[406]), .c ({signal_967, signal_146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_543 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_957, signal_548}), .a ({signal_956, signal_547}), .clk (clk), .r (Fresh[407]), .c ({signal_968, signal_145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_544 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_959, signal_550}), .a ({signal_958, signal_549}), .clk (clk), .r (Fresh[408]), .c ({signal_969, signal_144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(0)) cell_545 ( .s ({X_s1[7], X_s0[7]}), .b ({signal_961, signal_552}), .a ({signal_960, signal_551}), .clk (clk), .r (Fresh[409]), .c ({signal_970, signal_143}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_0 ( .clk (signal_1390), .D ({signal_970, signal_143}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1 ( .clk (signal_1390), .D ({signal_969, signal_144}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_2 ( .clk (signal_1390), .D ({signal_968, signal_145}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3 ( .clk (signal_1390), .D ({signal_967, signal_146}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_4 ( .clk (signal_1390), .D ({signal_966, signal_147}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_5 ( .clk (signal_1390), .D ({signal_965, signal_148}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_6 ( .clk (signal_1390), .D ({signal_964, signal_149}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_7 ( .clk (signal_1390), .D ({signal_963, signal_150}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
