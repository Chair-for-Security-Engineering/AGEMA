/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 16 time(s)  */

module sbox_HPC2_BDDsylvan_ClockGating_d4 (SI_s0, clk, SI_s1, SI_s2, SI_s3, SI_s4, Fresh, rst, SO_s0, SO_s1, SO_s2, SO_s3, SO_s4, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [7:0] SI_s4 ;
    input rst ;
    input [4099:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    output [7:0] SO_s4 ;
    output Synch ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_7149 ;

    /* cells in depth 0 */
    ClockGatingController #(17) cell_1337 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_7149 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_927 ( .s ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_928 ( .s ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_929 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_930 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_931 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_1375, signal_1374, signal_1373, signal_1372, signal_946}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_932 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_933 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_934 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_935 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_936 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_937 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_938 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_939 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_940 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_941 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_1415, signal_1414, signal_1413, signal_1412, signal_956}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_942 ( .s ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_943 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_1423, signal_1422, signal_1421, signal_1420, signal_958}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_944 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .c ({signal_1427, signal_1426, signal_1425, signal_1424, signal_959}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_945 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_1431, signal_1430, signal_1429, signal_1428, signal_960}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_946 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .c ({signal_1435, signal_1434, signal_1433, signal_1432, signal_961}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_947 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({signal_1439, signal_1438, signal_1437, signal_1436, signal_962}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_948 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_1443, signal_1442, signal_1441, signal_1440, signal_963}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_949 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({signal_1447, signal_1446, signal_1445, signal_1444, signal_964}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_950 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .c ({signal_1451, signal_1450, signal_1449, signal_1448, signal_965}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_951 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_1455, signal_1454, signal_1453, signal_1452, signal_966}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_952 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .c ({signal_1459, signal_1458, signal_1457, signal_1456, signal_967}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_953 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({signal_1463, signal_1462, signal_1461, signal_1460, signal_968}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_954 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_1467, signal_1466, signal_1465, signal_1464, signal_969}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_955 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({signal_1471, signal_1470, signal_1469, signal_1468, signal_970}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_956 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .c ({signal_1475, signal_1474, signal_1473, signal_1472, signal_971}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_957 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_1479, signal_1478, signal_1477, signal_1476, signal_972}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_958 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .c ({signal_1483, signal_1482, signal_1481, signal_1480, signal_973}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_959 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({signal_1487, signal_1486, signal_1485, signal_1484, signal_974}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_960 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_1491, signal_1490, signal_1489, signal_1488, signal_975}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_961 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({signal_1495, signal_1494, signal_1493, signal_1492, signal_976}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_962 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .c ({signal_1499, signal_1498, signal_1497, signal_1496, signal_977}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_963 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_964 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .c ({signal_1507, signal_1506, signal_1505, signal_1504, signal_979}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_965 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({signal_1511, signal_1510, signal_1509, signal_1508, signal_980}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_966 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_1515, signal_1514, signal_1513, signal_1512, signal_981}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_967 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .c ({signal_1519, signal_1518, signal_1517, signal_1516, signal_982}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_968 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .c ({signal_1523, signal_1522, signal_1521, signal_1520, signal_983}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_969 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_1527, signal_1526, signal_1525, signal_1524, signal_984}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_970 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .c ({signal_1531, signal_1530, signal_1529, signal_1528, signal_985}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_971 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .c ({signal_1535, signal_1534, signal_1533, signal_1532, signal_986}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_972 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_1539, signal_1538, signal_1537, signal_1536, signal_987}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_973 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .c ({signal_1543, signal_1542, signal_1541, signal_1540, signal_988}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_974 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .c ({signal_1547, signal_1546, signal_1545, signal_1544, signal_989}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_975 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_1551, signal_1550, signal_1549, signal_1548, signal_990}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_976 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .c ({signal_1555, signal_1554, signal_1553, signal_1552, signal_991}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_977 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .c ({signal_1559, signal_1558, signal_1557, signal_1556, signal_992}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_978 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_1563, signal_1562, signal_1561, signal_1560, signal_993}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_979 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .c ({signal_1567, signal_1566, signal_1565, signal_1564, signal_994}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_980 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .c ({signal_1571, signal_1570, signal_1569, signal_1568, signal_995}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_981 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_1575, signal_1574, signal_1573, signal_1572, signal_996}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_982 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .c ({signal_1579, signal_1578, signal_1577, signal_1576, signal_997}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_983 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .c ({signal_1583, signal_1582, signal_1581, signal_1580, signal_998}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_984 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_1587, signal_1586, signal_1585, signal_1584, signal_999}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_985 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .c ({signal_1591, signal_1590, signal_1589, signal_1588, signal_1000}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_986 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .c ({signal_1595, signal_1594, signal_1593, signal_1592, signal_1001}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_987 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_1599, signal_1598, signal_1597, signal_1596, signal_1002}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_988 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .c ({signal_1603, signal_1602, signal_1601, signal_1600, signal_1003}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_989 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .c ({signal_1607, signal_1606, signal_1605, signal_1604, signal_1004}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_990 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_1611, signal_1610, signal_1609, signal_1608, signal_1005}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_991 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .c ({signal_1615, signal_1614, signal_1613, signal_1612, signal_1006}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_992 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .c ({signal_1619, signal_1618, signal_1617, signal_1616, signal_1007}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_993 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_1623, signal_1622, signal_1621, signal_1620, signal_1008}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_994 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .c ({signal_1627, signal_1626, signal_1625, signal_1624, signal_1009}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_995 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .c ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_996 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_1635, signal_1634, signal_1633, signal_1632, signal_1011}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_997 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .c ({signal_1639, signal_1638, signal_1637, signal_1636, signal_1012}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_998 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .c ({signal_1643, signal_1642, signal_1641, signal_1640, signal_1013}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_999 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_1647, signal_1646, signal_1645, signal_1644, signal_1014}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1000 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .c ({signal_1651, signal_1650, signal_1649, signal_1648, signal_1015}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1001 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .c ({signal_1655, signal_1654, signal_1653, signal_1652, signal_1016}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1002 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_1659, signal_1658, signal_1657, signal_1656, signal_1017}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1003 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .c ({signal_1663, signal_1662, signal_1661, signal_1660, signal_1018}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1004 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .c ({signal_1667, signal_1666, signal_1665, signal_1664, signal_1019}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1005 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_1671, signal_1670, signal_1669, signal_1668, signal_1020}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1006 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .c ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1007 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .c ({signal_1679, signal_1678, signal_1677, signal_1676, signal_1022}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1008 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_1683, signal_1682, signal_1681, signal_1680, signal_1023}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1009 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .c ({signal_1687, signal_1686, signal_1685, signal_1684, signal_1024}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1010 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .c ({signal_1691, signal_1690, signal_1689, signal_1688, signal_1025}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1011 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_1695, signal_1694, signal_1693, signal_1692, signal_1026}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1012 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .c ({signal_1699, signal_1698, signal_1697, signal_1696, signal_1027}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1013 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .c ({signal_1703, signal_1702, signal_1701, signal_1700, signal_1028}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1014 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1707, signal_1706, signal_1705, signal_1704, signal_1029}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1015 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .c ({signal_1711, signal_1710, signal_1709, signal_1708, signal_1030}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1016 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890]}), .c ({signal_1715, signal_1714, signal_1713, signal_1712, signal_1031}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1017 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1719, signal_1718, signal_1717, signal_1716, signal_1032}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1018 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910]}), .c ({signal_1723, signal_1722, signal_1721, signal_1720, signal_1033}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1019 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .c ({signal_1727, signal_1726, signal_1725, signal_1724, signal_1034}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1020 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1731, signal_1730, signal_1729, signal_1728, signal_1035}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1021 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .c ({signal_1735, signal_1734, signal_1733, signal_1732, signal_1036}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1022 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950]}), .c ({signal_1739, signal_1738, signal_1737, signal_1736, signal_1037}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1023 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1743, signal_1742, signal_1741, signal_1740, signal_1038}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1024 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970]}), .c ({signal_1747, signal_1746, signal_1745, signal_1744, signal_1039}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1025 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .c ({signal_1751, signal_1750, signal_1749, signal_1748, signal_1040}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1026 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_1755, signal_1754, signal_1753, signal_1752, signal_1041}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1027 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .c ({signal_1759, signal_1758, signal_1757, signal_1756, signal_1042}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1028 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010]}), .c ({signal_1763, signal_1762, signal_1761, signal_1760, signal_1043}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1029 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_1767, signal_1766, signal_1765, signal_1764, signal_1044}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1030 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030]}), .c ({signal_1771, signal_1770, signal_1769, signal_1768, signal_1045}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1031 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .c ({signal_1775, signal_1774, signal_1773, signal_1772, signal_1046}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1032 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_1779, signal_1778, signal_1777, signal_1776, signal_1047}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1033 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .c ({signal_1783, signal_1782, signal_1781, signal_1780, signal_1048}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1034 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070]}), .c ({signal_1787, signal_1786, signal_1785, signal_1784, signal_1049}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1035 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1791, signal_1790, signal_1789, signal_1788, signal_1050}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1036 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090]}), .c ({signal_1795, signal_1794, signal_1793, signal_1792, signal_1051}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1037 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .c ({signal_1799, signal_1798, signal_1797, signal_1796, signal_1052}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1038 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1803, signal_1802, signal_1801, signal_1800, signal_1053}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1039 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .c ({signal_1807, signal_1806, signal_1805, signal_1804, signal_1054}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1040 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130]}), .c ({signal_1811, signal_1810, signal_1809, signal_1808, signal_1055}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1041 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1815, signal_1814, signal_1813, signal_1812, signal_1056}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1042 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150]}), .c ({signal_1819, signal_1818, signal_1817, signal_1816, signal_1057}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1043 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .c ({signal_1823, signal_1822, signal_1821, signal_1820, signal_1058}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1044 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1827, signal_1826, signal_1825, signal_1824, signal_1059}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1045 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .c ({signal_1831, signal_1830, signal_1829, signal_1828, signal_1060}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1046 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190]}), .c ({signal_1835, signal_1834, signal_1833, signal_1832, signal_1061}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1047 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1839, signal_1838, signal_1837, signal_1836, signal_1062}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1048 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210]}), .c ({signal_1843, signal_1842, signal_1841, signal_1840, signal_1063}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1049 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .c ({signal_1847, signal_1846, signal_1845, signal_1844, signal_1064}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1050 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_1851, signal_1850, signal_1849, signal_1848, signal_1065}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1051 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .clk ( clk ), .r ({Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .c ({signal_1855, signal_1854, signal_1853, signal_1852, signal_1066}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1052 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250]}), .c ({signal_1859, signal_1858, signal_1857, signal_1856, signal_1067}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1053 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1054 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270]}), .c ({signal_1867, signal_1866, signal_1865, signal_1864, signal_1069}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1055 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .c ({signal_1871, signal_1870, signal_1869, signal_1868, signal_1070}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1056 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_1875, signal_1874, signal_1873, signal_1872, signal_1071}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1057 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .c ({signal_1879, signal_1878, signal_1877, signal_1876, signal_1072}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1058 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310]}), .c ({signal_1883, signal_1882, signal_1881, signal_1880, signal_1073}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1059 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_1887, signal_1886, signal_1885, signal_1884, signal_1074}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1060 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330]}), .c ({signal_1891, signal_1890, signal_1889, signal_1888, signal_1075}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1061 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .c ({signal_1895, signal_1894, signal_1893, signal_1892, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1062 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_1899, signal_1898, signal_1897, signal_1896, signal_1077}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1063 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .c ({signal_1903, signal_1902, signal_1901, signal_1900, signal_1078}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1064 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370]}), .c ({signal_1907, signal_1906, signal_1905, signal_1904, signal_1079}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1065 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_1911, signal_1910, signal_1909, signal_1908, signal_1080}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1066 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390]}), .c ({signal_1915, signal_1914, signal_1913, signal_1912, signal_1081}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1067 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .c ({signal_1919, signal_1918, signal_1917, signal_1916, signal_1082}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1068 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_1923, signal_1922, signal_1921, signal_1920, signal_1083}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1069 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .c ({signal_1927, signal_1926, signal_1925, signal_1924, signal_1084}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1070 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430]}), .c ({signal_1931, signal_1930, signal_1929, signal_1928, signal_1085}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1071 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .clk ( clk ), .r ({Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_1935, signal_1934, signal_1933, signal_1932, signal_1086}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1072 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450]}), .c ({signal_1939, signal_1938, signal_1937, signal_1936, signal_1087}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1073 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .c ({signal_1943, signal_1942, signal_1941, signal_1940, signal_1088}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1074 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_1947, signal_1946, signal_1945, signal_1944, signal_1089}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1075 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .c ({signal_1951, signal_1950, signal_1949, signal_1948, signal_1090}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1076 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1351, signal_1350, signal_1349, signal_1348, signal_942}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490]}), .c ({signal_1955, signal_1954, signal_1953, signal_1952, signal_1091}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1077 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .clk ( clk ), .r ({Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_1959, signal_1958, signal_1957, signal_1956, signal_1092}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1078 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510]}), .c ({signal_1963, signal_1962, signal_1961, signal_1960, signal_1093}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1079 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .c ({signal_1967, signal_1966, signal_1965, signal_1964, signal_1094}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1080 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_1971, signal_1970, signal_1969, signal_1968, signal_1095}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1081 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({signal_1387, signal_1386, signal_1385, signal_1384, signal_949}), .clk ( clk ), .r ({Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .c ({signal_1975, signal_1974, signal_1973, signal_1972, signal_1096}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1082 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1383, signal_1382, signal_1381, signal_1380, signal_948}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550]}), .c ({signal_1979, signal_1978, signal_1977, signal_1976, signal_1097}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1083 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1399, signal_1398, signal_1397, signal_1396, signal_952}), .a ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .clk ( clk ), .r ({Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_1983, signal_1982, signal_1981, signal_1980, signal_1098}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1084 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1395, signal_1394, signal_1393, signal_1392, signal_951}), .a ({signal_1403, signal_1402, signal_1401, signal_1400, signal_953}), .clk ( clk ), .r ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570]}), .c ({signal_1987, signal_1986, signal_1985, signal_1984, signal_1099}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1085 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .c ({signal_1991, signal_1990, signal_1989, signal_1988, signal_1100}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1086 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1419, signal_1418, signal_1417, signal_1416, signal_957}), .clk ( clk ), .r ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_1995, signal_1994, signal_1993, signal_1992, signal_1101}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1087 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .a ({signal_1475, signal_1474, signal_1473, signal_1472, signal_971}), .clk ( clk ), .r ({Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .c ({signal_2003, signal_2002, signal_2001, signal_2000, signal_1102}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1088 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610]}), .c ({signal_2007, signal_2006, signal_2005, signal_2004, signal_1103}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1089 ( .s ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1411, signal_1410, signal_1409, signal_1408, signal_955}), .clk ( clk ), .r ({Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_2011, signal_2010, signal_2009, signal_2008, signal_1104}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1090 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1483, signal_1482, signal_1481, signal_1480, signal_973}), .a ({signal_1479, signal_1478, signal_1477, signal_1476, signal_972}), .clk ( clk ), .r ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630]}), .c ({signal_2015, signal_2014, signal_2013, signal_2012, signal_1105}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1091 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1491, signal_1490, signal_1489, signal_1488, signal_975}), .a ({signal_1487, signal_1486, signal_1485, signal_1484, signal_974}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .c ({signal_2019, signal_2018, signal_2017, signal_2016, signal_1106}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1092 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1499, signal_1498, signal_1497, signal_1496, signal_977}), .a ({signal_1495, signal_1494, signal_1493, signal_1492, signal_976}), .clk ( clk ), .r ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_2023, signal_2022, signal_2021, signal_2020, signal_1107}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1093 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1507, signal_1506, signal_1505, signal_1504, signal_979}), .a ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}), .clk ( clk ), .r ({Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .c ({signal_2027, signal_2026, signal_2025, signal_2024, signal_1108}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1094 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1515, signal_1514, signal_1513, signal_1512, signal_981}), .a ({signal_1511, signal_1510, signal_1509, signal_1508, signal_980}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670]}), .c ({signal_2031, signal_2030, signal_2029, signal_2028, signal_1109}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1095 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1511, signal_1510, signal_1509, signal_1508, signal_980}), .a ({signal_1519, signal_1518, signal_1517, signal_1516, signal_982}), .clk ( clk ), .r ({Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_2035, signal_2034, signal_2033, signal_2032, signal_1110}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1096 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1523, signal_1522, signal_1521, signal_1520, signal_983}), .a ({signal_1415, signal_1414, signal_1413, signal_1412, signal_956}), .clk ( clk ), .r ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690]}), .c ({signal_2039, signal_2038, signal_2037, signal_2036, signal_1111}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1097 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1531, signal_1530, signal_1529, signal_1528, signal_985}), .a ({signal_1527, signal_1526, signal_1525, signal_1524, signal_984}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .c ({signal_2043, signal_2042, signal_2041, signal_2040, signal_1112}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1098 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1539, signal_1538, signal_1537, signal_1536, signal_987}), .a ({signal_1535, signal_1534, signal_1533, signal_1532, signal_986}), .clk ( clk ), .r ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_2047, signal_2046, signal_2045, signal_2044, signal_1113}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1099 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1423, signal_1422, signal_1421, signal_1420, signal_958}), .a ({signal_1543, signal_1542, signal_1541, signal_1540, signal_988}), .clk ( clk ), .r ({Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .c ({signal_2051, signal_2050, signal_2049, signal_2048, signal_1114}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1100 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1551, signal_1550, signal_1549, signal_1548, signal_990}), .a ({signal_1547, signal_1546, signal_1545, signal_1544, signal_989}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730]}), .c ({signal_2055, signal_2054, signal_2053, signal_2052, signal_1115}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1101 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1555, signal_1554, signal_1553, signal_1552, signal_991}), .a ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}), .clk ( clk ), .r ({Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_2059, signal_2058, signal_2057, signal_2056, signal_1116}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1102 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1563, signal_1562, signal_1561, signal_1560, signal_993}), .a ({signal_1559, signal_1558, signal_1557, signal_1556, signal_992}), .clk ( clk ), .r ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750]}), .c ({signal_2063, signal_2062, signal_2061, signal_2060, signal_1117}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1103 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1571, signal_1570, signal_1569, signal_1568, signal_995}), .a ({signal_1567, signal_1566, signal_1565, signal_1564, signal_994}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .c ({signal_2067, signal_2066, signal_2065, signal_2064, signal_1118}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1104 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1579, signal_1578, signal_1577, signal_1576, signal_997}), .a ({signal_1575, signal_1574, signal_1573, signal_1572, signal_996}), .clk ( clk ), .r ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_2071, signal_2070, signal_2069, signal_2068, signal_1119}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1105 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1587, signal_1586, signal_1585, signal_1584, signal_999}), .a ({signal_1583, signal_1582, signal_1581, signal_1580, signal_998}), .clk ( clk ), .r ({Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .c ({signal_2075, signal_2074, signal_2073, signal_2072, signal_1120}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1106 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1595, signal_1594, signal_1593, signal_1592, signal_1001}), .a ({signal_1591, signal_1590, signal_1589, signal_1588, signal_1000}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790]}), .c ({signal_2079, signal_2078, signal_2077, signal_2076, signal_1121}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1107 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1603, signal_1602, signal_1601, signal_1600, signal_1003}), .a ({signal_1599, signal_1598, signal_1597, signal_1596, signal_1002}), .clk ( clk ), .r ({Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_2083, signal_2082, signal_2081, signal_2080, signal_1122}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1108 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1527, signal_1526, signal_1525, signal_1524, signal_984}), .a ({signal_1607, signal_1606, signal_1605, signal_1604, signal_1004}), .clk ( clk ), .r ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810]}), .c ({signal_2087, signal_2086, signal_2085, signal_2084, signal_1123}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1109 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1615, signal_1614, signal_1613, signal_1612, signal_1006}), .a ({signal_1611, signal_1610, signal_1609, signal_1608, signal_1005}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .c ({signal_2091, signal_2090, signal_2089, signal_2088, signal_1124}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1110 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1623, signal_1622, signal_1621, signal_1620, signal_1008}), .a ({signal_1619, signal_1618, signal_1617, signal_1616, signal_1007}), .clk ( clk ), .r ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_2095, signal_2094, signal_2093, signal_2092, signal_1125}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1111 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}), .a ({signal_1627, signal_1626, signal_1625, signal_1624, signal_1009}), .clk ( clk ), .r ({Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .c ({signal_2099, signal_2098, signal_2097, signal_2096, signal_1126}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1112 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1635, signal_1634, signal_1633, signal_1632, signal_1011}), .a ({signal_1427, signal_1426, signal_1425, signal_1424, signal_959}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850]}), .c ({signal_2103, signal_2102, signal_2101, signal_2100, signal_1127}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1113 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1643, signal_1642, signal_1641, signal_1640, signal_1013}), .a ({signal_1639, signal_1638, signal_1637, signal_1636, signal_1012}), .clk ( clk ), .r ({Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_2107, signal_2106, signal_2105, signal_2104, signal_1128}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1114 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1651, signal_1650, signal_1649, signal_1648, signal_1015}), .a ({signal_1647, signal_1646, signal_1645, signal_1644, signal_1014}), .clk ( clk ), .r ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870]}), .c ({signal_2111, signal_2110, signal_2109, signal_2108, signal_1129}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1115 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1659, signal_1658, signal_1657, signal_1656, signal_1017}), .a ({signal_1655, signal_1654, signal_1653, signal_1652, signal_1016}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .c ({signal_2115, signal_2114, signal_2113, signal_2112, signal_1130}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1116 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1663, signal_1662, signal_1661, signal_1660, signal_1018}), .a ({signal_1599, signal_1598, signal_1597, signal_1596, signal_1002}), .clk ( clk ), .r ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_2119, signal_2118, signal_2117, signal_2116, signal_1131}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1117 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}), .a ({signal_1495, signal_1494, signal_1493, signal_1492, signal_976}), .clk ( clk ), .r ({Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .c ({signal_2123, signal_2122, signal_2121, signal_2120, signal_1132}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1118 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1671, signal_1670, signal_1669, signal_1668, signal_1020}), .a ({signal_1667, signal_1666, signal_1665, signal_1664, signal_1019}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910]}), .c ({signal_2127, signal_2126, signal_2125, signal_2124, signal_1133}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1119 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .clk ( clk ), .r ({Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_2131, signal_2130, signal_2129, signal_2128, signal_1134}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1120 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1431, signal_1430, signal_1429, signal_1428, signal_960}), .a ({signal_1655, signal_1654, signal_1653, signal_1652, signal_1016}), .clk ( clk ), .r ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930]}), .c ({signal_2135, signal_2134, signal_2133, signal_2132, signal_1135}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1121 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}), .a ({signal_1435, signal_1434, signal_1433, signal_1432, signal_961}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .c ({signal_2139, signal_2138, signal_2137, signal_2136, signal_1136}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1122 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1491, signal_1490, signal_1489, signal_1488, signal_975}), .a ({signal_1439, signal_1438, signal_1437, signal_1436, signal_962}), .clk ( clk ), .r ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_2143, signal_2142, signal_2141, signal_2140, signal_1137}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1123 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1415, signal_1414, signal_1413, signal_1412, signal_956}), .a ({signal_1679, signal_1678, signal_1677, signal_1676, signal_1022}), .clk ( clk ), .r ({Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .c ({signal_2147, signal_2146, signal_2145, signal_2144, signal_1138}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1124 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1687, signal_1686, signal_1685, signal_1684, signal_1024}), .a ({signal_1683, signal_1682, signal_1681, signal_1680, signal_1023}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970]}), .c ({signal_2151, signal_2150, signal_2149, signal_2148, signal_1139}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1125 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1435, signal_1434, signal_1433, signal_1432, signal_961}), .a ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}), .clk ( clk ), .r ({Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_2155, signal_2154, signal_2153, signal_2152, signal_1140}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1126 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}), .a ({signal_1691, signal_1690, signal_1689, signal_1688, signal_1025}), .clk ( clk ), .r ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990]}), .c ({signal_2159, signal_2158, signal_2157, signal_2156, signal_1141}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1127 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1699, signal_1698, signal_1697, signal_1696, signal_1027}), .a ({signal_1695, signal_1694, signal_1693, signal_1692, signal_1026}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .c ({signal_2163, signal_2162, signal_2161, signal_2160, signal_1142}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1128 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1443, signal_1442, signal_1441, signal_1440, signal_963}), .a ({signal_1703, signal_1702, signal_1701, signal_1700, signal_1028}), .clk ( clk ), .r ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_2167, signal_2166, signal_2165, signal_2164, signal_1143}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1129 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1707, signal_1706, signal_1705, signal_1704, signal_1029}), .a ({signal_1447, signal_1446, signal_1445, signal_1444, signal_964}), .clk ( clk ), .r ({Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .c ({signal_2171, signal_2170, signal_2169, signal_2168, signal_1144}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1130 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1715, signal_1714, signal_1713, signal_1712, signal_1031}), .a ({signal_1711, signal_1710, signal_1709, signal_1708, signal_1030}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030]}), .c ({signal_2175, signal_2174, signal_2173, signal_2172, signal_1145}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1131 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1723, signal_1722, signal_1721, signal_1720, signal_1033}), .a ({signal_1719, signal_1718, signal_1717, signal_1716, signal_1032}), .clk ( clk ), .r ({Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_2179, signal_2178, signal_2177, signal_2176, signal_1146}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1132 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1731, signal_1730, signal_1729, signal_1728, signal_1035}), .a ({signal_1727, signal_1726, signal_1725, signal_1724, signal_1034}), .clk ( clk ), .r ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050]}), .c ({signal_2183, signal_2182, signal_2181, signal_2180, signal_1147}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1133 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1499, signal_1498, signal_1497, signal_1496, signal_977}), .a ({signal_1735, signal_1734, signal_1733, signal_1732, signal_1036}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .c ({signal_2187, signal_2186, signal_2185, signal_2184, signal_1148}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1134 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1743, signal_1742, signal_1741, signal_1740, signal_1038}), .a ({signal_1739, signal_1738, signal_1737, signal_1736, signal_1037}), .clk ( clk ), .r ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_2191, signal_2190, signal_2189, signal_2188, signal_1149}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1135 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1707, signal_1706, signal_1705, signal_1704, signal_1029}), .a ({signal_1747, signal_1746, signal_1745, signal_1744, signal_1039}), .clk ( clk ), .r ({Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .c ({signal_2195, signal_2194, signal_2193, signal_2192, signal_1150}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1136 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1751, signal_1750, signal_1749, signal_1748, signal_1040}), .a ({signal_1703, signal_1702, signal_1701, signal_1700, signal_1028}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090]}), .c ({signal_2199, signal_2198, signal_2197, signal_2196, signal_1151}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1137 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1755, signal_1754, signal_1753, signal_1752, signal_1041}), .a ({signal_1643, signal_1642, signal_1641, signal_1640, signal_1013}), .clk ( clk ), .r ({Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_2203, signal_2202, signal_2201, signal_2200, signal_1152}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1138 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1759, signal_1758, signal_1757, signal_1756, signal_1042}), .a ({signal_1563, signal_1562, signal_1561, signal_1560, signal_993}), .clk ( clk ), .r ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110]}), .c ({signal_2207, signal_2206, signal_2205, signal_2204, signal_1153}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1139 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1767, signal_1766, signal_1765, signal_1764, signal_1044}), .a ({signal_1763, signal_1762, signal_1761, signal_1760, signal_1043}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .c ({signal_2211, signal_2210, signal_2209, signal_2208, signal_1154}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1140 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1771, signal_1770, signal_1769, signal_1768, signal_1045}), .a ({signal_1591, signal_1590, signal_1589, signal_1588, signal_1000}), .clk ( clk ), .r ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_2215, signal_2214, signal_2213, signal_2212, signal_1155}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1141 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1775, signal_1774, signal_1773, signal_1772, signal_1046}), .a ({signal_1707, signal_1706, signal_1705, signal_1704, signal_1029}), .clk ( clk ), .r ({Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .c ({signal_2219, signal_2218, signal_2217, signal_2216, signal_1156}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1142 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1783, signal_1782, signal_1781, signal_1780, signal_1048}), .a ({signal_1779, signal_1778, signal_1777, signal_1776, signal_1047}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150]}), .c ({signal_2223, signal_2222, signal_2221, signal_2220, signal_1157}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1143 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1791, signal_1790, signal_1789, signal_1788, signal_1050}), .a ({signal_1787, signal_1786, signal_1785, signal_1784, signal_1049}), .clk ( clk ), .r ({Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_2227, signal_2226, signal_2225, signal_2224, signal_1158}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1144 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1439, signal_1438, signal_1437, signal_1436, signal_962}), .a ({signal_1795, signal_1794, signal_1793, signal_1792, signal_1051}), .clk ( clk ), .r ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170]}), .c ({signal_2231, signal_2230, signal_2229, signal_2228, signal_1159}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1145 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1775, signal_1774, signal_1773, signal_1772, signal_1046}), .a ({signal_1579, signal_1578, signal_1577, signal_1576, signal_997}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .c ({signal_2235, signal_2234, signal_2233, signal_2232, signal_1160}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1146 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1535, signal_1534, signal_1533, signal_1532, signal_986}), .a ({signal_1799, signal_1798, signal_1797, signal_1796, signal_1052}), .clk ( clk ), .r ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_2239, signal_2238, signal_2237, signal_2236, signal_1161}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1147 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}), .a ({signal_1527, signal_1526, signal_1525, signal_1524, signal_984}), .clk ( clk ), .r ({Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .c ({signal_2243, signal_2242, signal_2241, signal_2240, signal_1162}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1148 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1715, signal_1714, signal_1713, signal_1712, signal_1031}), .a ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210]}), .c ({signal_2247, signal_2246, signal_2245, signal_2244, signal_1163}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1149 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}), .a ({signal_1803, signal_1802, signal_1801, signal_1800, signal_1053}), .clk ( clk ), .r ({Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_2251, signal_2250, signal_2249, signal_2248, signal_1164}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1150 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1807, signal_1806, signal_1805, signal_1804, signal_1054}), .a ({signal_1511, signal_1510, signal_1509, signal_1508, signal_980}), .clk ( clk ), .r ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230]}), .c ({signal_2255, signal_2254, signal_2253, signal_2252, signal_1165}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1151 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1723, signal_1722, signal_1721, signal_1720, signal_1033}), .a ({signal_1811, signal_1810, signal_1809, signal_1808, signal_1055}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .c ({signal_2259, signal_2258, signal_2257, signal_2256, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1152 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1819, signal_1818, signal_1817, signal_1816, signal_1057}), .a ({signal_1815, signal_1814, signal_1813, signal_1812, signal_1056}), .clk ( clk ), .r ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_2263, signal_2262, signal_2261, signal_2260, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1153 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1619, signal_1618, signal_1617, signal_1616, signal_1007}), .a ({signal_1823, signal_1822, signal_1821, signal_1820, signal_1058}), .clk ( clk ), .r ({Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .c ({signal_2267, signal_2266, signal_2265, signal_2264, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1154 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1511, signal_1510, signal_1509, signal_1508, signal_980}), .a ({signal_1827, signal_1826, signal_1825, signal_1824, signal_1059}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270]}), .c ({signal_2271, signal_2270, signal_2269, signal_2268, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1155 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1671, signal_1670, signal_1669, signal_1668, signal_1020}), .a ({signal_1451, signal_1450, signal_1449, signal_1448, signal_965}), .clk ( clk ), .r ({Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_2275, signal_2274, signal_2273, signal_2272, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1156 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1831, signal_1830, signal_1829, signal_1828, signal_1060}), .a ({signal_1687, signal_1686, signal_1685, signal_1684, signal_1024}), .clk ( clk ), .r ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290]}), .c ({signal_2279, signal_2278, signal_2277, signal_2276, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1157 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1431, signal_1430, signal_1429, signal_1428, signal_960}), .a ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .c ({signal_2283, signal_2282, signal_2281, signal_2280, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1158 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1499, signal_1498, signal_1497, signal_1496, signal_977}), .a ({signal_1835, signal_1834, signal_1833, signal_1832, signal_1061}), .clk ( clk ), .r ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_2287, signal_2286, signal_2285, signal_2284, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1159 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1639, signal_1638, signal_1637, signal_1636, signal_1012}), .a ({signal_1519, signal_1518, signal_1517, signal_1516, signal_982}), .clk ( clk ), .r ({Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .c ({signal_2291, signal_2290, signal_2289, signal_2288, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1160 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1751, signal_1750, signal_1749, signal_1748, signal_1040}), .a ({signal_1839, signal_1838, signal_1837, signal_1836, signal_1062}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330]}), .c ({signal_2295, signal_2294, signal_2293, signal_2292, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1161 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1643, signal_1642, signal_1641, signal_1640, signal_1013}), .a ({signal_1843, signal_1842, signal_1841, signal_1840, signal_1063}), .clk ( clk ), .r ({Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_2299, signal_2298, signal_2297, signal_2296, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1162 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1851, signal_1850, signal_1849, signal_1848, signal_1065}), .a ({signal_1847, signal_1846, signal_1845, signal_1844, signal_1064}), .clk ( clk ), .r ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350]}), .c ({signal_2303, signal_2302, signal_2301, signal_2300, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1163 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1855, signal_1854, signal_1853, signal_1852, signal_1066}), .a ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .c ({signal_2307, signal_2306, signal_2305, signal_2304, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1164 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1859, signal_1858, signal_1857, signal_1856, signal_1067}), .a ({signal_1655, signal_1654, signal_1653, signal_1652, signal_1016}), .clk ( clk ), .r ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_2311, signal_2310, signal_2309, signal_2308, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1165 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1823, signal_1822, signal_1821, signal_1820, signal_1058}), .a ({signal_1375, signal_1374, signal_1373, signal_1372, signal_946}), .clk ( clk ), .r ({Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .c ({signal_2315, signal_2314, signal_2313, signal_2312, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1166 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1867, signal_1866, signal_1865, signal_1864, signal_1069}), .a ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390]}), .c ({signal_2319, signal_2318, signal_2317, signal_2316, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1167 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .a ({signal_1871, signal_1870, signal_1869, signal_1868, signal_1070}), .clk ( clk ), .r ({Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_2323, signal_2322, signal_2321, signal_2320, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1168 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1875, signal_1874, signal_1873, signal_1872, signal_1071}), .a ({signal_1803, signal_1802, signal_1801, signal_1800, signal_1053}), .clk ( clk ), .r ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410]}), .c ({signal_2327, signal_2326, signal_2325, signal_2324, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1169 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1483, signal_1482, signal_1481, signal_1480, signal_973}), .a ({signal_1559, signal_1558, signal_1557, signal_1556, signal_992}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .c ({signal_2331, signal_2330, signal_2329, signal_2328, signal_1184}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1170 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1519, signal_1518, signal_1517, signal_1516, signal_982}), .a ({signal_1879, signal_1878, signal_1877, signal_1876, signal_1072}), .clk ( clk ), .r ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_2335, signal_2334, signal_2333, signal_2332, signal_1185}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1171 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1555, signal_1554, signal_1553, signal_1552, signal_991}), .a ({signal_1751, signal_1750, signal_1749, signal_1748, signal_1040}), .clk ( clk ), .r ({Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .c ({signal_2339, signal_2338, signal_2337, signal_2336, signal_1186}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1172 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1479, signal_1478, signal_1477, signal_1476, signal_972}), .a ({signal_1627, signal_1626, signal_1625, signal_1624, signal_1009}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450]}), .c ({signal_2343, signal_2342, signal_2341, signal_2340, signal_1187}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1173 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1495, signal_1494, signal_1493, signal_1492, signal_976}), .a ({signal_1799, signal_1798, signal_1797, signal_1796, signal_1052}), .clk ( clk ), .r ({Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_2347, signal_2346, signal_2345, signal_2344, signal_1188}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1174 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1883, signal_1882, signal_1881, signal_1880, signal_1073}), .a ({signal_1675, signal_1674, signal_1673, signal_1672, signal_1021}), .clk ( clk ), .r ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470]}), .c ({signal_2351, signal_2350, signal_2349, signal_2348, signal_1189}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1175 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1831, signal_1830, signal_1829, signal_1828, signal_1060}), .a ({signal_1367, signal_1366, signal_1365, signal_1364, signal_945}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .c ({signal_2355, signal_2354, signal_2353, signal_2352, signal_1190}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1176 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1887, signal_1886, signal_1885, signal_1884, signal_1074}), .a ({signal_1523, signal_1522, signal_1521, signal_1520, signal_983}), .clk ( clk ), .r ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_2359, signal_2358, signal_2357, signal_2356, signal_1191}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1177 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1895, signal_1894, signal_1893, signal_1892, signal_1076}), .a ({signal_1891, signal_1890, signal_1889, signal_1888, signal_1075}), .clk ( clk ), .r ({Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .c ({signal_2363, signal_2362, signal_2361, signal_2360, signal_1192}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1178 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}), .a ({signal_1899, signal_1898, signal_1897, signal_1896, signal_1077}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510]}), .c ({signal_2367, signal_2366, signal_2365, signal_2364, signal_1193}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1179 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1563, signal_1562, signal_1561, signal_1560, signal_993}), .a ({signal_1355, signal_1354, signal_1353, signal_1352, signal_943}), .clk ( clk ), .r ({Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_2371, signal_2370, signal_2369, signal_2368, signal_1194}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1180 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1907, signal_1906, signal_1905, signal_1904, signal_1079}), .a ({signal_1903, signal_1902, signal_1901, signal_1900, signal_1078}), .clk ( clk ), .r ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530]}), .c ({signal_2375, signal_2374, signal_2373, signal_2372, signal_1195}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1181 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1727, signal_1726, signal_1725, signal_1724, signal_1034}), .a ({signal_1503, signal_1502, signal_1501, signal_1500, signal_978}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .c ({signal_2379, signal_2378, signal_2377, signal_2376, signal_1196}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1182 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1507, signal_1506, signal_1505, signal_1504, signal_979}), .a ({signal_1911, signal_1910, signal_1909, signal_1908, signal_1080}), .clk ( clk ), .r ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_2383, signal_2382, signal_2381, signal_2380, signal_1197}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1183 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1667, signal_1666, signal_1665, signal_1664, signal_1019}), .a ({signal_1455, signal_1454, signal_1453, signal_1452, signal_966}), .clk ( clk ), .r ({Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .c ({signal_2387, signal_2386, signal_2385, signal_2384, signal_1198}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1184 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1919, signal_1918, signal_1917, signal_1916, signal_1082}), .a ({signal_1915, signal_1914, signal_1913, signal_1912, signal_1081}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570]}), .c ({signal_2391, signal_2390, signal_2389, signal_2388, signal_1199}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1185 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1923, signal_1922, signal_1921, signal_1920, signal_1083}), .a ({signal_1391, signal_1390, signal_1389, signal_1388, signal_950}), .clk ( clk ), .r ({Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_2395, signal_2394, signal_2393, signal_2392, signal_1200}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1186 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1699, signal_1698, signal_1697, signal_1696, signal_1027}), .a ({signal_1927, signal_1926, signal_1925, signal_1924, signal_1084}), .clk ( clk ), .r ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590]}), .c ({signal_2399, signal_2398, signal_2397, signal_2396, signal_1201}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1187 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1363, signal_1362, signal_1361, signal_1360, signal_944}), .a ({signal_1875, signal_1874, signal_1873, signal_1872, signal_1071}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .c ({signal_2403, signal_2402, signal_2401, signal_2400, signal_1202}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1188 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1931, signal_1930, signal_1929, signal_1928, signal_1085}), .a ({signal_1799, signal_1798, signal_1797, signal_1796, signal_1052}), .clk ( clk ), .r ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_2407, signal_2406, signal_2405, signal_2404, signal_1203}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1189 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1939, signal_1938, signal_1937, signal_1936, signal_1087}), .a ({signal_1935, signal_1934, signal_1933, signal_1932, signal_1086}), .clk ( clk ), .r ({Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .c ({signal_2411, signal_2410, signal_2409, signal_2408, signal_1204}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1190 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1899, signal_1898, signal_1897, signal_1896, signal_1077}), .a ({signal_1447, signal_1446, signal_1445, signal_1444, signal_964}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630]}), .c ({signal_2415, signal_2414, signal_2413, signal_2412, signal_1205}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1191 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1943, signal_1942, signal_1941, signal_1940, signal_1088}), .a ({signal_1551, signal_1550, signal_1549, signal_1548, signal_990}), .clk ( clk ), .r ({Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_2419, signal_2418, signal_2417, signal_2416, signal_1206}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1192 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1903, signal_1902, signal_1901, signal_1900, signal_1078}), .a ({signal_1947, signal_1946, signal_1945, signal_1944, signal_1089}), .clk ( clk ), .r ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650]}), .c ({signal_2423, signal_2422, signal_2421, signal_2420, signal_1207}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1193 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1931, signal_1930, signal_1929, signal_1928, signal_1085}), .a ({signal_1531, signal_1530, signal_1529, signal_1528, signal_985}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .c ({signal_2427, signal_2426, signal_2425, signal_2424, signal_1208}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1194 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1955, signal_1954, signal_1953, signal_1952, signal_1091}), .a ({signal_1951, signal_1950, signal_1949, signal_1948, signal_1090}), .clk ( clk ), .r ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_2431, signal_2430, signal_2429, signal_2428, signal_1209}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1195 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1703, signal_1702, signal_1701, signal_1700, signal_1028}), .a ({signal_1775, signal_1774, signal_1773, signal_1772, signal_1046}), .clk ( clk ), .r ({Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .c ({signal_2435, signal_2434, signal_2433, signal_2432, signal_1210}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1196 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1539, signal_1538, signal_1537, signal_1536, signal_987}), .a ({signal_1427, signal_1426, signal_1425, signal_1424, signal_959}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690]}), .c ({signal_2439, signal_2438, signal_2437, signal_2436, signal_1211}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1197 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1959, signal_1958, signal_1957, signal_1956, signal_1092}), .a ({signal_1799, signal_1798, signal_1797, signal_1796, signal_1052}), .clk ( clk ), .r ({Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_2443, signal_2442, signal_2441, signal_2440, signal_1212}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1198 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1459, signal_1458, signal_1457, signal_1456, signal_967}), .a ({signal_1919, signal_1918, signal_1917, signal_1916, signal_1082}), .clk ( clk ), .r ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710]}), .c ({signal_2447, signal_2446, signal_2445, signal_2444, signal_1213}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1199 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}), .a ({signal_1463, signal_1462, signal_1461, signal_1460, signal_968}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .c ({signal_2451, signal_2450, signal_2449, signal_2448, signal_1214}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1200 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1963, signal_1962, signal_1961, signal_1960, signal_1093}), .a ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}), .clk ( clk ), .r ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_2455, signal_2454, signal_2453, signal_2452, signal_1215}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1201 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_1643, signal_1642, signal_1641, signal_1640, signal_1013}), .clk ( clk ), .r ({Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .c ({signal_2459, signal_2458, signal_2457, signal_2456, signal_1216}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1202 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1967, signal_1966, signal_1965, signal_1964, signal_1094}), .a ({signal_1803, signal_1802, signal_1801, signal_1800, signal_1053}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750]}), .c ({signal_2463, signal_2462, signal_2461, signal_2460, signal_1217}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1203 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1971, signal_1970, signal_1969, signal_1968, signal_1095}), .a ({signal_1759, signal_1758, signal_1757, signal_1756, signal_1042}), .clk ( clk ), .r ({Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_2467, signal_2466, signal_2465, signal_2464, signal_1218}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1204 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1379, signal_1378, signal_1377, signal_1376, signal_947}), .a ({signal_1875, signal_1874, signal_1873, signal_1872, signal_1071}), .clk ( clk ), .r ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770]}), .c ({signal_2471, signal_2470, signal_2469, signal_2468, signal_1219}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1205 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1975, signal_1974, signal_1973, signal_1972, signal_1096}), .a ({signal_1859, signal_1858, signal_1857, signal_1856, signal_1067}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .c ({signal_2475, signal_2474, signal_2473, signal_2472, signal_1220}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1206 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1947, signal_1946, signal_1945, signal_1944, signal_1089}), .a ({signal_1655, signal_1654, signal_1653, signal_1652, signal_1016}), .clk ( clk ), .r ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_2479, signal_2478, signal_2477, signal_2476, signal_1221}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1207 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1979, signal_1978, signal_1977, signal_1976, signal_1097}), .a ({signal_1407, signal_1406, signal_1405, signal_1404, signal_954}), .clk ( clk ), .r ({Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .c ({signal_2483, signal_2482, signal_2481, signal_2480, signal_1222}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1208 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1467, signal_1466, signal_1465, signal_1464, signal_969}), .a ({signal_1983, signal_1982, signal_1981, signal_1980, signal_1098}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810]}), .c ({signal_2487, signal_2486, signal_2485, signal_2484, signal_1223}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1209 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1987, signal_1986, signal_1985, signal_1984, signal_1099}), .a ({signal_1471, signal_1470, signal_1469, signal_1468, signal_970}), .clk ( clk ), .r ({Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_2491, signal_2490, signal_2489, signal_2488, signal_1224}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1210 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1991, signal_1990, signal_1989, signal_1988, signal_1100}), .a ({signal_1971, signal_1970, signal_1969, signal_1968, signal_1095}), .clk ( clk ), .r ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830]}), .c ({signal_2495, signal_2494, signal_2493, signal_2492, signal_1225}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1211 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1995, signal_1994, signal_1993, signal_1992, signal_1101}), .a ({signal_1863, signal_1862, signal_1861, signal_1860, signal_1068}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .c ({signal_2499, signal_2498, signal_2497, signal_2496, signal_1226}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1212 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1619, signal_1618, signal_1617, signal_1616, signal_1007}), .a ({signal_1639, signal_1638, signal_1637, signal_1636, signal_1012}), .clk ( clk ), .r ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_2503, signal_2502, signal_2501, signal_2500, signal_1227}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1213 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1939, signal_1938, signal_1937, signal_1936, signal_1087}), .a ({signal_1439, signal_1438, signal_1437, signal_1436, signal_962}), .clk ( clk ), .r ({Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .c ({signal_2507, signal_2506, signal_2505, signal_2504, signal_1228}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1214 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2007, signal_2006, signal_2005, signal_2004, signal_1103}), .a ({signal_1631, signal_1630, signal_1629, signal_1628, signal_1010}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870]}), .c ({signal_2511, signal_2510, signal_2509, signal_2508, signal_1229}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1215 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1599, signal_1598, signal_1597, signal_1596, signal_1002}), .a ({signal_2011, signal_2010, signal_2009, signal_2008, signal_1104}), .clk ( clk ), .r ({Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_2515, signal_2514, signal_2513, signal_2512, signal_1230}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1216 ( .s ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_1807, signal_1806, signal_1805, signal_1804, signal_1054}), .a ({signal_1595, signal_1594, signal_1593, signal_1592, signal_1001}), .clk ( clk ), .r ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890]}), .c ({signal_2519, signal_2518, signal_2517, signal_2516, signal_1231}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1217 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2019, signal_2018, signal_2017, signal_2016, signal_1106}), .a ({signal_2015, signal_2014, signal_2013, signal_2012, signal_1105}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .c ({signal_2527, signal_2526, signal_2525, signal_2524, signal_1232}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1218 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2027, signal_2026, signal_2025, signal_2024, signal_1108}), .a ({signal_2023, signal_2022, signal_2021, signal_2020, signal_1107}), .clk ( clk ), .r ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_2531, signal_2530, signal_2529, signal_2528, signal_1233}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1219 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2035, signal_2034, signal_2033, signal_2032, signal_1110}), .a ({signal_2031, signal_2030, signal_2029, signal_2028, signal_1109}), .clk ( clk ), .r ({Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .c ({signal_2535, signal_2534, signal_2533, signal_2532, signal_1234}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1220 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2043, signal_2042, signal_2041, signal_2040, signal_1112}), .a ({signal_2039, signal_2038, signal_2037, signal_2036, signal_1111}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930]}), .c ({signal_2539, signal_2538, signal_2537, signal_2536, signal_1235}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1221 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2051, signal_2050, signal_2049, signal_2048, signal_1114}), .a ({signal_2047, signal_2046, signal_2045, signal_2044, signal_1113}), .clk ( clk ), .r ({Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_2543, signal_2542, signal_2541, signal_2540, signal_1236}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1222 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2059, signal_2058, signal_2057, signal_2056, signal_1116}), .a ({signal_2055, signal_2054, signal_2053, signal_2052, signal_1115}), .clk ( clk ), .r ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950]}), .c ({signal_2547, signal_2546, signal_2545, signal_2544, signal_1237}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1223 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2067, signal_2066, signal_2065, signal_2064, signal_1118}), .a ({signal_2063, signal_2062, signal_2061, signal_2060, signal_1117}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .c ({signal_2551, signal_2550, signal_2549, signal_2548, signal_1238}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1224 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2075, signal_2074, signal_2073, signal_2072, signal_1120}), .a ({signal_2071, signal_2070, signal_2069, signal_2068, signal_1119}), .clk ( clk ), .r ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_2555, signal_2554, signal_2553, signal_2552, signal_1239}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1225 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2083, signal_2082, signal_2081, signal_2080, signal_1122}), .a ({signal_2079, signal_2078, signal_2077, signal_2076, signal_1121}), .clk ( clk ), .r ({Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .c ({signal_2559, signal_2558, signal_2557, signal_2556, signal_1240}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1226 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2091, signal_2090, signal_2089, signal_2088, signal_1124}), .a ({signal_2087, signal_2086, signal_2085, signal_2084, signal_1123}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990]}), .c ({signal_2563, signal_2562, signal_2561, signal_2560, signal_1241}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1227 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2099, signal_2098, signal_2097, signal_2096, signal_1126}), .a ({signal_2095, signal_2094, signal_2093, signal_2092, signal_1125}), .clk ( clk ), .r ({Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_2567, signal_2566, signal_2565, signal_2564, signal_1242}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1228 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2107, signal_2106, signal_2105, signal_2104, signal_1128}), .a ({signal_2103, signal_2102, signal_2101, signal_2100, signal_1127}), .clk ( clk ), .r ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010]}), .c ({signal_2571, signal_2570, signal_2569, signal_2568, signal_1243}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1229 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2115, signal_2114, signal_2113, signal_2112, signal_1130}), .a ({signal_2111, signal_2110, signal_2109, signal_2108, signal_1129}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .c ({signal_2575, signal_2574, signal_2573, signal_2572, signal_1244}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1230 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2123, signal_2122, signal_2121, signal_2120, signal_1132}), .a ({signal_2119, signal_2118, signal_2117, signal_2116, signal_1131}), .clk ( clk ), .r ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_2579, signal_2578, signal_2577, signal_2576, signal_1245}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1231 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2131, signal_2130, signal_2129, signal_2128, signal_1134}), .a ({signal_2127, signal_2126, signal_2125, signal_2124, signal_1133}), .clk ( clk ), .r ({Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .c ({signal_2583, signal_2582, signal_2581, signal_2580, signal_1246}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1232 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2139, signal_2138, signal_2137, signal_2136, signal_1136}), .a ({signal_2135, signal_2134, signal_2133, signal_2132, signal_1135}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050]}), .c ({signal_2587, signal_2586, signal_2585, signal_2584, signal_1247}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1233 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2147, signal_2146, signal_2145, signal_2144, signal_1138}), .a ({signal_2143, signal_2142, signal_2141, signal_2140, signal_1137}), .clk ( clk ), .r ({Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_2591, signal_2590, signal_2589, signal_2588, signal_1248}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1234 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2155, signal_2154, signal_2153, signal_2152, signal_1140}), .a ({signal_2151, signal_2150, signal_2149, signal_2148, signal_1139}), .clk ( clk ), .r ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070]}), .c ({signal_2595, signal_2594, signal_2593, signal_2592, signal_1249}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1235 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2163, signal_2162, signal_2161, signal_2160, signal_1142}), .a ({signal_2159, signal_2158, signal_2157, signal_2156, signal_1141}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .c ({signal_2599, signal_2598, signal_2597, signal_2596, signal_1250}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1236 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2171, signal_2170, signal_2169, signal_2168, signal_1144}), .a ({signal_2167, signal_2166, signal_2165, signal_2164, signal_1143}), .clk ( clk ), .r ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_2603, signal_2602, signal_2601, signal_2600, signal_1251}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1237 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2179, signal_2178, signal_2177, signal_2176, signal_1146}), .a ({signal_2175, signal_2174, signal_2173, signal_2172, signal_1145}), .clk ( clk ), .r ({Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .c ({signal_2607, signal_2606, signal_2605, signal_2604, signal_1252}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1238 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2187, signal_2186, signal_2185, signal_2184, signal_1148}), .a ({signal_2183, signal_2182, signal_2181, signal_2180, signal_1147}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110]}), .c ({signal_2611, signal_2610, signal_2609, signal_2608, signal_1253}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1239 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2195, signal_2194, signal_2193, signal_2192, signal_1150}), .a ({signal_2191, signal_2190, signal_2189, signal_2188, signal_1149}), .clk ( clk ), .r ({Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_2615, signal_2614, signal_2613, signal_2612, signal_1254}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1240 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2203, signal_2202, signal_2201, signal_2200, signal_1152}), .a ({signal_2199, signal_2198, signal_2197, signal_2196, signal_1151}), .clk ( clk ), .r ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130]}), .c ({signal_2619, signal_2618, signal_2617, signal_2616, signal_1255}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1241 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2211, signal_2210, signal_2209, signal_2208, signal_1154}), .a ({signal_2207, signal_2206, signal_2205, signal_2204, signal_1153}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .c ({signal_2623, signal_2622, signal_2621, signal_2620, signal_1256}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1242 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2219, signal_2218, signal_2217, signal_2216, signal_1156}), .a ({signal_2215, signal_2214, signal_2213, signal_2212, signal_1155}), .clk ( clk ), .r ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_2627, signal_2626, signal_2625, signal_2624, signal_1257}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1243 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2227, signal_2226, signal_2225, signal_2224, signal_1158}), .a ({signal_2223, signal_2222, signal_2221, signal_2220, signal_1157}), .clk ( clk ), .r ({Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .c ({signal_2631, signal_2630, signal_2629, signal_2628, signal_1258}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1244 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2235, signal_2234, signal_2233, signal_2232, signal_1160}), .a ({signal_2231, signal_2230, signal_2229, signal_2228, signal_1159}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170]}), .c ({signal_2635, signal_2634, signal_2633, signal_2632, signal_1259}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1245 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2243, signal_2242, signal_2241, signal_2240, signal_1162}), .a ({signal_2239, signal_2238, signal_2237, signal_2236, signal_1161}), .clk ( clk ), .r ({Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_2639, signal_2638, signal_2637, signal_2636, signal_1260}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1246 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2251, signal_2250, signal_2249, signal_2248, signal_1164}), .a ({signal_2247, signal_2246, signal_2245, signal_2244, signal_1163}), .clk ( clk ), .r ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190]}), .c ({signal_2643, signal_2642, signal_2641, signal_2640, signal_1261}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1247 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2259, signal_2258, signal_2257, signal_2256, signal_1166}), .a ({signal_2255, signal_2254, signal_2253, signal_2252, signal_1165}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .c ({signal_2647, signal_2646, signal_2645, signal_2644, signal_1262}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1248 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2267, signal_2266, signal_2265, signal_2264, signal_1168}), .a ({signal_2263, signal_2262, signal_2261, signal_2260, signal_1167}), .clk ( clk ), .r ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_2651, signal_2650, signal_2649, signal_2648, signal_1263}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1249 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2275, signal_2274, signal_2273, signal_2272, signal_1170}), .a ({signal_2271, signal_2270, signal_2269, signal_2268, signal_1169}), .clk ( clk ), .r ({Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .c ({signal_2655, signal_2654, signal_2653, signal_2652, signal_1264}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1250 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2283, signal_2282, signal_2281, signal_2280, signal_1172}), .a ({signal_2279, signal_2278, signal_2277, signal_2276, signal_1171}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230]}), .c ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1265}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1251 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2291, signal_2290, signal_2289, signal_2288, signal_1174}), .a ({signal_2287, signal_2286, signal_2285, signal_2284, signal_1173}), .clk ( clk ), .r ({Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1266}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1252 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2299, signal_2298, signal_2297, signal_2296, signal_1176}), .a ({signal_2295, signal_2294, signal_2293, signal_2292, signal_1175}), .clk ( clk ), .r ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250]}), .c ({signal_2667, signal_2666, signal_2665, signal_2664, signal_1267}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1253 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2307, signal_2306, signal_2305, signal_2304, signal_1178}), .a ({signal_2303, signal_2302, signal_2301, signal_2300, signal_1177}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .c ({signal_2671, signal_2670, signal_2669, signal_2668, signal_1268}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1254 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2315, signal_2314, signal_2313, signal_2312, signal_1180}), .a ({signal_2311, signal_2310, signal_2309, signal_2308, signal_1179}), .clk ( clk ), .r ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1269}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1255 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2323, signal_2322, signal_2321, signal_2320, signal_1182}), .a ({signal_2319, signal_2318, signal_2317, signal_2316, signal_1181}), .clk ( clk ), .r ({Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .c ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1270}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1256 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2331, signal_2330, signal_2329, signal_2328, signal_1184}), .a ({signal_2327, signal_2326, signal_2325, signal_2324, signal_1183}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290]}), .c ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1271}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1257 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2339, signal_2338, signal_2337, signal_2336, signal_1186}), .a ({signal_2335, signal_2334, signal_2333, signal_2332, signal_1185}), .clk ( clk ), .r ({Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1272}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1258 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2347, signal_2346, signal_2345, signal_2344, signal_1188}), .a ({signal_2343, signal_2342, signal_2341, signal_2340, signal_1187}), .clk ( clk ), .r ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310]}), .c ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1273}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1259 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2355, signal_2354, signal_2353, signal_2352, signal_1190}), .a ({signal_2351, signal_2350, signal_2349, signal_2348, signal_1189}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .c ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1274}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1260 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2363, signal_2362, signal_2361, signal_2360, signal_1192}), .a ({signal_2359, signal_2358, signal_2357, signal_2356, signal_1191}), .clk ( clk ), .r ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1275}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1261 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2371, signal_2370, signal_2369, signal_2368, signal_1194}), .a ({signal_2367, signal_2366, signal_2365, signal_2364, signal_1193}), .clk ( clk ), .r ({Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .c ({signal_2703, signal_2702, signal_2701, signal_2700, signal_1276}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1262 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2379, signal_2378, signal_2377, signal_2376, signal_1196}), .a ({signal_2375, signal_2374, signal_2373, signal_2372, signal_1195}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350]}), .c ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1277}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1263 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2387, signal_2386, signal_2385, signal_2384, signal_1198}), .a ({signal_2383, signal_2382, signal_2381, signal_2380, signal_1197}), .clk ( clk ), .r ({Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_2711, signal_2710, signal_2709, signal_2708, signal_1278}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1264 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2395, signal_2394, signal_2393, signal_2392, signal_1200}), .a ({signal_2391, signal_2390, signal_2389, signal_2388, signal_1199}), .clk ( clk ), .r ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370]}), .c ({signal_2715, signal_2714, signal_2713, signal_2712, signal_1279}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1265 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2403, signal_2402, signal_2401, signal_2400, signal_1202}), .a ({signal_2399, signal_2398, signal_2397, signal_2396, signal_1201}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .c ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1280}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1266 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2411, signal_2410, signal_2409, signal_2408, signal_1204}), .a ({signal_2407, signal_2406, signal_2405, signal_2404, signal_1203}), .clk ( clk ), .r ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1281}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1267 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2419, signal_2418, signal_2417, signal_2416, signal_1206}), .a ({signal_2415, signal_2414, signal_2413, signal_2412, signal_1205}), .clk ( clk ), .r ({Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .c ({signal_2727, signal_2726, signal_2725, signal_2724, signal_1282}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1268 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2427, signal_2426, signal_2425, signal_2424, signal_1208}), .a ({signal_2423, signal_2422, signal_2421, signal_2420, signal_1207}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410]}), .c ({signal_2731, signal_2730, signal_2729, signal_2728, signal_1283}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1269 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2435, signal_2434, signal_2433, signal_2432, signal_1210}), .a ({signal_2431, signal_2430, signal_2429, signal_2428, signal_1209}), .clk ( clk ), .r ({Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_2735, signal_2734, signal_2733, signal_2732, signal_1284}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1270 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2443, signal_2442, signal_2441, signal_2440, signal_1212}), .a ({signal_2439, signal_2438, signal_2437, signal_2436, signal_1211}), .clk ( clk ), .r ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430]}), .c ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1285}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1271 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2451, signal_2450, signal_2449, signal_2448, signal_1214}), .a ({signal_2447, signal_2446, signal_2445, signal_2444, signal_1213}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .c ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1286}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1272 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2459, signal_2458, signal_2457, signal_2456, signal_1216}), .a ({signal_2455, signal_2454, signal_2453, signal_2452, signal_1215}), .clk ( clk ), .r ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_2747, signal_2746, signal_2745, signal_2744, signal_1287}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1273 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2467, signal_2466, signal_2465, signal_2464, signal_1218}), .a ({signal_2463, signal_2462, signal_2461, signal_2460, signal_1217}), .clk ( clk ), .r ({Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .c ({signal_2751, signal_2750, signal_2749, signal_2748, signal_1288}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1274 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2475, signal_2474, signal_2473, signal_2472, signal_1220}), .a ({signal_2471, signal_2470, signal_2469, signal_2468, signal_1219}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470]}), .c ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1289}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1275 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2483, signal_2482, signal_2481, signal_2480, signal_1222}), .a ({signal_2479, signal_2478, signal_2477, signal_2476, signal_1221}), .clk ( clk ), .r ({Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_2759, signal_2758, signal_2757, signal_2756, signal_1290}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1276 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2491, signal_2490, signal_2489, signal_2488, signal_1224}), .a ({signal_2487, signal_2486, signal_2485, signal_2484, signal_1223}), .clk ( clk ), .r ({Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490]}), .c ({signal_2763, signal_2762, signal_2761, signal_2760, signal_1291}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1277 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2499, signal_2498, signal_2497, signal_2496, signal_1226}), .a ({signal_2495, signal_2494, signal_2493, signal_2492, signal_1225}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500]}), .c ({signal_2767, signal_2766, signal_2765, signal_2764, signal_1292}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1278 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2507, signal_2506, signal_2505, signal_2504, signal_1228}), .a ({signal_2503, signal_2502, signal_2501, signal_2500, signal_1227}), .clk ( clk ), .r ({Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_2771, signal_2770, signal_2769, signal_2768, signal_1293}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1279 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2511, signal_2510, signal_2509, signal_2508, signal_1229}), .a ({signal_2003, signal_2002, signal_2001, signal_2000, signal_1102}), .clk ( clk ), .r ({Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520]}), .c ({signal_2775, signal_2774, signal_2773, signal_2772, signal_1294}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1280 ( .s ({SI_s4[4], SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2519, signal_2518, signal_2517, signal_2516, signal_1231}), .a ({signal_2515, signal_2514, signal_2513, signal_2512, signal_1230}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530]}), .c ({signal_2779, signal_2778, signal_2777, signal_2776, signal_1295}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1281 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2531, signal_2530, signal_2529, signal_2528, signal_1233}), .a ({signal_2527, signal_2526, signal_2525, signal_2524, signal_1232}), .clk ( clk ), .r ({Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_2787, signal_2786, signal_2785, signal_2784, signal_1296}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1282 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2539, signal_2538, signal_2537, signal_2536, signal_1235}), .a ({signal_2535, signal_2534, signal_2533, signal_2532, signal_1234}), .clk ( clk ), .r ({Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550]}), .c ({signal_2791, signal_2790, signal_2789, signal_2788, signal_1297}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1283 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2547, signal_2546, signal_2545, signal_2544, signal_1237}), .a ({signal_2543, signal_2542, signal_2541, signal_2540, signal_1236}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560]}), .c ({signal_2795, signal_2794, signal_2793, signal_2792, signal_1298}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1284 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2555, signal_2554, signal_2553, signal_2552, signal_1239}), .a ({signal_2551, signal_2550, signal_2549, signal_2548, signal_1238}), .clk ( clk ), .r ({Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_2799, signal_2798, signal_2797, signal_2796, signal_1299}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1285 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2563, signal_2562, signal_2561, signal_2560, signal_1241}), .a ({signal_2559, signal_2558, signal_2557, signal_2556, signal_1240}), .clk ( clk ), .r ({Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580]}), .c ({signal_2803, signal_2802, signal_2801, signal_2800, signal_1300}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1286 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2571, signal_2570, signal_2569, signal_2568, signal_1243}), .a ({signal_2567, signal_2566, signal_2565, signal_2564, signal_1242}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590]}), .c ({signal_2807, signal_2806, signal_2805, signal_2804, signal_1301}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1287 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2579, signal_2578, signal_2577, signal_2576, signal_1245}), .a ({signal_2575, signal_2574, signal_2573, signal_2572, signal_1244}), .clk ( clk ), .r ({Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_2811, signal_2810, signal_2809, signal_2808, signal_1302}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1288 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2587, signal_2586, signal_2585, signal_2584, signal_1247}), .a ({signal_2583, signal_2582, signal_2581, signal_2580, signal_1246}), .clk ( clk ), .r ({Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610]}), .c ({signal_2815, signal_2814, signal_2813, signal_2812, signal_1303}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1289 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2595, signal_2594, signal_2593, signal_2592, signal_1249}), .a ({signal_2591, signal_2590, signal_2589, signal_2588, signal_1248}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620]}), .c ({signal_2819, signal_2818, signal_2817, signal_2816, signal_1304}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1290 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2603, signal_2602, signal_2601, signal_2600, signal_1251}), .a ({signal_2599, signal_2598, signal_2597, signal_2596, signal_1250}), .clk ( clk ), .r ({Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_2823, signal_2822, signal_2821, signal_2820, signal_1305}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1291 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2611, signal_2610, signal_2609, signal_2608, signal_1253}), .a ({signal_2607, signal_2606, signal_2605, signal_2604, signal_1252}), .clk ( clk ), .r ({Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640]}), .c ({signal_2827, signal_2826, signal_2825, signal_2824, signal_1306}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1292 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2619, signal_2618, signal_2617, signal_2616, signal_1255}), .a ({signal_2615, signal_2614, signal_2613, signal_2612, signal_1254}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650]}), .c ({signal_2831, signal_2830, signal_2829, signal_2828, signal_1307}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1293 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2627, signal_2626, signal_2625, signal_2624, signal_1257}), .a ({signal_2623, signal_2622, signal_2621, signal_2620, signal_1256}), .clk ( clk ), .r ({Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_2835, signal_2834, signal_2833, signal_2832, signal_1308}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1294 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2635, signal_2634, signal_2633, signal_2632, signal_1259}), .a ({signal_2631, signal_2630, signal_2629, signal_2628, signal_1258}), .clk ( clk ), .r ({Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670]}), .c ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1309}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1295 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2643, signal_2642, signal_2641, signal_2640, signal_1261}), .a ({signal_2639, signal_2638, signal_2637, signal_2636, signal_1260}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680]}), .c ({signal_2843, signal_2842, signal_2841, signal_2840, signal_1310}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1296 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2651, signal_2650, signal_2649, signal_2648, signal_1263}), .a ({signal_2647, signal_2646, signal_2645, signal_2644, signal_1262}), .clk ( clk ), .r ({Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_2847, signal_2846, signal_2845, signal_2844, signal_1311}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1297 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2659, signal_2658, signal_2657, signal_2656, signal_1265}), .a ({signal_2655, signal_2654, signal_2653, signal_2652, signal_1264}), .clk ( clk ), .r ({Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700]}), .c ({signal_2851, signal_2850, signal_2849, signal_2848, signal_1312}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1298 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2667, signal_2666, signal_2665, signal_2664, signal_1267}), .a ({signal_2663, signal_2662, signal_2661, signal_2660, signal_1266}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710]}), .c ({signal_2855, signal_2854, signal_2853, signal_2852, signal_1313}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1299 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2675, signal_2674, signal_2673, signal_2672, signal_1269}), .a ({signal_2671, signal_2670, signal_2669, signal_2668, signal_1268}), .clk ( clk ), .r ({Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_2859, signal_2858, signal_2857, signal_2856, signal_1314}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1300 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2683, signal_2682, signal_2681, signal_2680, signal_1271}), .a ({signal_2679, signal_2678, signal_2677, signal_2676, signal_1270}), .clk ( clk ), .r ({Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730]}), .c ({signal_2863, signal_2862, signal_2861, signal_2860, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1301 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2691, signal_2690, signal_2689, signal_2688, signal_1273}), .a ({signal_2687, signal_2686, signal_2685, signal_2684, signal_1272}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740]}), .c ({signal_2867, signal_2866, signal_2865, signal_2864, signal_1316}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1302 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2699, signal_2698, signal_2697, signal_2696, signal_1275}), .a ({signal_2695, signal_2694, signal_2693, signal_2692, signal_1274}), .clk ( clk ), .r ({Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_2871, signal_2870, signal_2869, signal_2868, signal_1317}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1303 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2707, signal_2706, signal_2705, signal_2704, signal_1277}), .a ({signal_2703, signal_2702, signal_2701, signal_2700, signal_1276}), .clk ( clk ), .r ({Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760]}), .c ({signal_2875, signal_2874, signal_2873, signal_2872, signal_1318}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1304 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2715, signal_2714, signal_2713, signal_2712, signal_1279}), .a ({signal_2711, signal_2710, signal_2709, signal_2708, signal_1278}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770]}), .c ({signal_2879, signal_2878, signal_2877, signal_2876, signal_1319}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1305 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2723, signal_2722, signal_2721, signal_2720, signal_1281}), .a ({signal_2719, signal_2718, signal_2717, signal_2716, signal_1280}), .clk ( clk ), .r ({Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_2883, signal_2882, signal_2881, signal_2880, signal_1320}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1306 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2731, signal_2730, signal_2729, signal_2728, signal_1283}), .a ({signal_2727, signal_2726, signal_2725, signal_2724, signal_1282}), .clk ( clk ), .r ({Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790]}), .c ({signal_2887, signal_2886, signal_2885, signal_2884, signal_1321}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1307 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2739, signal_2738, signal_2737, signal_2736, signal_1285}), .a ({signal_2735, signal_2734, signal_2733, signal_2732, signal_1284}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800]}), .c ({signal_2891, signal_2890, signal_2889, signal_2888, signal_1322}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1308 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2747, signal_2746, signal_2745, signal_2744, signal_1287}), .a ({signal_2743, signal_2742, signal_2741, signal_2740, signal_1286}), .clk ( clk ), .r ({Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_2895, signal_2894, signal_2893, signal_2892, signal_1323}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1309 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2755, signal_2754, signal_2753, signal_2752, signal_1289}), .a ({signal_2751, signal_2750, signal_2749, signal_2748, signal_1288}), .clk ( clk ), .r ({Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820]}), .c ({signal_2899, signal_2898, signal_2897, signal_2896, signal_1324}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1310 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2763, signal_2762, signal_2761, signal_2760, signal_1291}), .a ({signal_2759, signal_2758, signal_2757, signal_2756, signal_1290}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830]}), .c ({signal_2903, signal_2902, signal_2901, signal_2900, signal_1325}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1311 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2771, signal_2770, signal_2769, signal_2768, signal_1293}), .a ({signal_2767, signal_2766, signal_2765, signal_2764, signal_1292}), .clk ( clk ), .r ({Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_2907, signal_2906, signal_2905, signal_2904, signal_1326}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1312 ( .s ({SI_s4[5], SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2779, signal_2778, signal_2777, signal_2776, signal_1295}), .a ({signal_2775, signal_2774, signal_2773, signal_2772, signal_1294}), .clk ( clk ), .r ({Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850]}), .c ({signal_2911, signal_2910, signal_2909, signal_2908, signal_1327}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1313 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2791, signal_2790, signal_2789, signal_2788, signal_1297}), .a ({signal_2787, signal_2786, signal_2785, signal_2784, signal_1296}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860]}), .c ({signal_2919, signal_2918, signal_2917, signal_2916, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1314 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2799, signal_2798, signal_2797, signal_2796, signal_1299}), .a ({signal_2795, signal_2794, signal_2793, signal_2792, signal_1298}), .clk ( clk ), .r ({Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_2923, signal_2922, signal_2921, signal_2920, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1315 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2807, signal_2806, signal_2805, signal_2804, signal_1301}), .a ({signal_2803, signal_2802, signal_2801, signal_2800, signal_1300}), .clk ( clk ), .r ({Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880]}), .c ({signal_2927, signal_2926, signal_2925, signal_2924, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1316 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2815, signal_2814, signal_2813, signal_2812, signal_1303}), .a ({signal_2811, signal_2810, signal_2809, signal_2808, signal_1302}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890]}), .c ({signal_2931, signal_2930, signal_2929, signal_2928, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1317 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2823, signal_2822, signal_2821, signal_2820, signal_1305}), .a ({signal_2819, signal_2818, signal_2817, signal_2816, signal_1304}), .clk ( clk ), .r ({Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_2935, signal_2934, signal_2933, signal_2932, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1318 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2831, signal_2830, signal_2829, signal_2828, signal_1307}), .a ({signal_2827, signal_2826, signal_2825, signal_2824, signal_1306}), .clk ( clk ), .r ({Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910]}), .c ({signal_2939, signal_2938, signal_2937, signal_2936, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1319 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2839, signal_2838, signal_2837, signal_2836, signal_1309}), .a ({signal_2835, signal_2834, signal_2833, signal_2832, signal_1308}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920]}), .c ({signal_2943, signal_2942, signal_2941, signal_2940, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1320 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2847, signal_2846, signal_2845, signal_2844, signal_1311}), .a ({signal_2843, signal_2842, signal_2841, signal_2840, signal_1310}), .clk ( clk ), .r ({Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_2947, signal_2946, signal_2945, signal_2944, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1321 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2855, signal_2854, signal_2853, signal_2852, signal_1313}), .a ({signal_2851, signal_2850, signal_2849, signal_2848, signal_1312}), .clk ( clk ), .r ({Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940]}), .c ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1322 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2863, signal_2862, signal_2861, signal_2860, signal_1315}), .a ({signal_2859, signal_2858, signal_2857, signal_2856, signal_1314}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950]}), .c ({signal_2955, signal_2954, signal_2953, signal_2952, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1323 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2871, signal_2870, signal_2869, signal_2868, signal_1317}), .a ({signal_2867, signal_2866, signal_2865, signal_2864, signal_1316}), .clk ( clk ), .r ({Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1324 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2879, signal_2878, signal_2877, signal_2876, signal_1319}), .a ({signal_2875, signal_2874, signal_2873, signal_2872, signal_1318}), .clk ( clk ), .r ({Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970]}), .c ({signal_2963, signal_2962, signal_2961, signal_2960, signal_1339}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1325 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2887, signal_2886, signal_2885, signal_2884, signal_1321}), .a ({signal_2883, signal_2882, signal_2881, signal_2880, signal_1320}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980]}), .c ({signal_2967, signal_2966, signal_2965, signal_2964, signal_1340}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1326 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2895, signal_2894, signal_2893, signal_2892, signal_1323}), .a ({signal_2891, signal_2890, signal_2889, signal_2888, signal_1322}), .clk ( clk ), .r ({Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1341}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1327 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2903, signal_2902, signal_2901, signal_2900, signal_1325}), .a ({signal_2899, signal_2898, signal_2897, signal_2896, signal_1324}), .clk ( clk ), .r ({Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000]}), .c ({signal_2975, signal_2974, signal_2973, signal_2972, signal_1342}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1328 ( .s ({SI_s4[6], SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2911, signal_2910, signal_2909, signal_2908, signal_1327}), .a ({signal_2907, signal_2906, signal_2905, signal_2904, signal_1326}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010]}), .c ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1343}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1329 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2923, signal_2922, signal_2921, signal_2920, signal_1329}), .a ({signal_2919, signal_2918, signal_2917, signal_2916, signal_1328}), .clk ( clk ), .r ({Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_2987, signal_2986, signal_2985, signal_2984, signal_30}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1330 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2931, signal_2930, signal_2929, signal_2928, signal_1331}), .a ({signal_2927, signal_2926, signal_2925, signal_2924, signal_1330}), .clk ( clk ), .r ({Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030]}), .c ({signal_2991, signal_2990, signal_2989, signal_2988, signal_29}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1331 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2939, signal_2938, signal_2937, signal_2936, signal_1333}), .a ({signal_2935, signal_2934, signal_2933, signal_2932, signal_1332}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040]}), .c ({signal_2995, signal_2994, signal_2993, signal_2992, signal_28}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1332 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2947, signal_2946, signal_2945, signal_2944, signal_1335}), .a ({signal_2943, signal_2942, signal_2941, signal_2940, signal_1334}), .clk ( clk ), .r ({Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_2999, signal_2998, signal_2997, signal_2996, signal_27}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1333 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2955, signal_2954, signal_2953, signal_2952, signal_1337}), .a ({signal_2951, signal_2950, signal_2949, signal_2948, signal_1336}), .clk ( clk ), .r ({Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060]}), .c ({signal_3003, signal_3002, signal_3001, signal_3000, signal_26}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1334 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2963, signal_2962, signal_2961, signal_2960, signal_1339}), .a ({signal_2959, signal_2958, signal_2957, signal_2956, signal_1338}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070]}), .c ({signal_3007, signal_3006, signal_3005, signal_3004, signal_25}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1335 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2971, signal_2970, signal_2969, signal_2968, signal_1341}), .a ({signal_2967, signal_2966, signal_2965, signal_2964, signal_1340}), .clk ( clk ), .r ({Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_3011, signal_3010, signal_3009, signal_3008, signal_24}) ) ;
    mux2_HPC2 #(.security_order(4), .pipeline(0)) cell_1336 ( .s ({SI_s4[7], SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2979, signal_2978, signal_2977, signal_2976, signal_1343}), .a ({signal_2975, signal_2974, signal_2973, signal_2972, signal_1342}), .clk ( clk ), .r ({Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090]}), .c ({signal_3015, signal_3014, signal_3013, signal_3012, signal_23}) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(0)) cell_0 ( .clk ( signal_7149 ), .D ({signal_3015, signal_3014, signal_3013, signal_3012, signal_23}), .Q ({SO_s4[7], SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_1 ( .clk ( signal_7149 ), .D ({signal_3011, signal_3010, signal_3009, signal_3008, signal_24}), .Q ({SO_s4[6], SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_2 ( .clk ( signal_7149 ), .D ({signal_3007, signal_3006, signal_3005, signal_3004, signal_25}), .Q ({SO_s4[5], SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_3 ( .clk ( signal_7149 ), .D ({signal_3003, signal_3002, signal_3001, signal_3000, signal_26}), .Q ({SO_s4[4], SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_4 ( .clk ( signal_7149 ), .D ({signal_2999, signal_2998, signal_2997, signal_2996, signal_27}), .Q ({SO_s4[3], SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_5 ( .clk ( signal_7149 ), .D ({signal_2995, signal_2994, signal_2993, signal_2992, signal_28}), .Q ({SO_s4[2], SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_6 ( .clk ( signal_7149 ), .D ({signal_2991, signal_2990, signal_2989, signal_2988, signal_29}), .Q ({SO_s4[1], SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(0)) cell_7 ( .clk ( signal_7149 ), .D ({signal_2987, signal_2986, signal_2985, signal_2984, signal_30}), .Q ({SO_s4[0], SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
