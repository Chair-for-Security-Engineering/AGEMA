/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 34 time(s)  */

module sbox_HPC2_AIG_ClockGating_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, rst, SO_s0, SO_s1, SO_s2, SO_s3, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input rst ;
    input [5273:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    output Synch ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_12089 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(0)) cell_927 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2397, signal_2396, signal_2395, signal_942}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_928 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2403, signal_2402, signal_2401, signal_943}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_929 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_930 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_931 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_932 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_933 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_934 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) cell_949 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .c ({signal_2484, signal_2483, signal_2482, signal_964}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) cell_950 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .c ({signal_2487, signal_2486, signal_2485, signal_965}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_962 ( .a ({signal_2484, signal_2483, signal_2482, signal_964}), .b ({signal_2523, signal_2522, signal_2521, signal_977}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_963 ( .a ({signal_2487, signal_2486, signal_2485, signal_965}), .b ({signal_2526, signal_2525, signal_2524, signal_978}) ) ;
    ClockGatingController #(35) cell_2385 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_12089 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_935 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_2442, signal_2441, signal_2440, signal_950}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_936 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_2445, signal_2444, signal_2443, signal_951}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_937 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_2448, signal_2447, signal_2446, signal_952}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_938 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_2451, signal_2450, signal_2449, signal_953}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_939 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_2454, signal_2453, signal_2452, signal_954}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_940 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_2457, signal_2456, signal_2455, signal_955}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_941 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_2460, signal_2459, signal_2458, signal_956}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_942 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_2463, signal_2462, signal_2461, signal_957}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_943 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_2466, signal_2465, signal_2464, signal_958}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_944 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_2469, signal_2468, signal_2467, signal_959}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_945 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_2472, signal_2471, signal_2470, signal_960}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_946 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_2475, signal_2474, signal_2473, signal_961}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_947 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_2478, signal_2477, signal_2476, signal_962}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_948 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_2481, signal_2480, signal_2479, signal_963}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_951 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2490, signal_2489, signal_2488, signal_966}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_952 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2493, signal_2492, signal_2491, signal_967}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_953 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2496, signal_2495, signal_2494, signal_968}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_954 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2499, signal_2498, signal_2497, signal_969}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_955 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2502, signal_2501, signal_2500, signal_970}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_956 ( .a ({signal_2460, signal_2459, signal_2458, signal_956}), .b ({signal_2505, signal_2504, signal_2503, signal_971}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_957 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2508, signal_2507, signal_2506, signal_972}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_958 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2511, signal_2510, signal_2509, signal_973}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_959 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2514, signal_2513, signal_2512, signal_974}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_960 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2517, signal_2516, signal_2515, signal_975}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_961 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2520, signal_2519, signal_2518, signal_976}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_964 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_2529, signal_2528, signal_2527, signal_979}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_965 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_2532, signal_2531, signal_2530, signal_980}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_966 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_2535, signal_2534, signal_2533, signal_981}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_967 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_2538, signal_2537, signal_2536, signal_982}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_968 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_2541, signal_2540, signal_2539, signal_983}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_969 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2403, signal_2402, signal_2401, signal_943}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_2544, signal_2543, signal_2542, signal_984}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_970 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_2547, signal_2546, signal_2545, signal_985}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_971 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_2550, signal_2549, signal_2548, signal_986}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_972 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_2553, signal_2552, signal_2551, signal_987}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_973 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_2556, signal_2555, signal_2554, signal_988}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_974 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_2559, signal_2558, signal_2557, signal_989}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_975 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_2562, signal_2561, signal_2560, signal_990}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_976 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_2565, signal_2564, signal_2563, signal_991}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_977 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_2568, signal_2567, signal_2566, signal_992}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_978 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_2571, signal_2570, signal_2569, signal_993}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_979 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_2574, signal_2573, signal_2572, signal_994}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_980 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_2577, signal_2576, signal_2575, signal_995}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_981 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_2580, signal_2579, signal_2578, signal_996}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_982 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_2583, signal_2582, signal_2581, signal_997}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_983 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_2586, signal_2585, signal_2584, signal_998}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_984 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_2589, signal_2588, signal_2587, signal_999}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_985 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_2592, signal_2591, signal_2590, signal_1000}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_986 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2403, signal_2402, signal_2401, signal_943}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_2595, signal_2594, signal_2593, signal_1001}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_987 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_2598, signal_2597, signal_2596, signal_1002}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_989 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_2604, signal_2603, signal_2602, signal_1004}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_990 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_2607, signal_2606, signal_2605, signal_1005}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_991 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_2610, signal_2609, signal_2608, signal_1006}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_992 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_2613, signal_2612, signal_2611, signal_1007}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_993 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_2616, signal_2615, signal_2614, signal_1008}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_994 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_2619, signal_2618, signal_2617, signal_1009}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_995 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_2622, signal_2621, signal_2620, signal_1010}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_996 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_2625, signal_2624, signal_2623, signal_1011}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_997 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_2628, signal_2627, signal_2626, signal_1012}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_998 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_2631, signal_2630, signal_2629, signal_1013}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1000 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_2637, signal_2636, signal_2635, signal_1015}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1001 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_2640, signal_2639, signal_2638, signal_1016}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1002 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_2643, signal_2642, signal_2641, signal_1017}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1003 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_2646, signal_2645, signal_2644, signal_1018}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1016 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2685, signal_2684, signal_2683, signal_1031}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1017 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2688, signal_2687, signal_2686, signal_1032}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1018 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2691, signal_2690, signal_2689, signal_1033}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1019 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2694, signal_2693, signal_2692, signal_1034}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1020 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2697, signal_2696, signal_2695, signal_1035}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1021 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_2700, signal_2699, signal_2698, signal_1036}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1022 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2703, signal_2702, signal_2701, signal_1037}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1023 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2706, signal_2705, signal_2704, signal_1038}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1024 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2709, signal_2708, signal_2707, signal_1039}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1025 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2712, signal_2711, signal_2710, signal_1040}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1026 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2715, signal_2714, signal_2713, signal_1041}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1027 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2718, signal_2717, signal_2716, signal_1042}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1028 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1029 ( .a ({signal_2580, signal_2579, signal_2578, signal_996}), .b ({signal_2724, signal_2723, signal_2722, signal_1044}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1030 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1031 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1032 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2733, signal_2732, signal_2731, signal_1047}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1034 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2739, signal_2738, signal_2737, signal_1049}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1035 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2742, signal_2741, signal_2740, signal_1050}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1036 ( .a ({signal_2610, signal_2609, signal_2608, signal_1006}), .b ({signal_2745, signal_2744, signal_2743, signal_1051}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1037 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1038 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1039 ( .a ({signal_2631, signal_2630, signal_2629, signal_1013}), .b ({signal_2754, signal_2753, signal_2752, signal_1054}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1041 ( .a ({signal_2637, signal_2636, signal_2635, signal_1015}), .b ({signal_2760, signal_2759, signal_2758, signal_1056}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1042 ( .a ({signal_2640, signal_2639, signal_2638, signal_1016}), .b ({signal_2763, signal_2762, signal_2761, signal_1057}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1043 ( .a ({signal_2643, signal_2642, signal_2641, signal_1017}), .b ({signal_2766, signal_2765, signal_2764, signal_1058}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_988 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_2601, signal_2600, signal_2599, signal_1003}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_999 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2457, signal_2456, signal_2455, signal_955}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_2634, signal_2633, signal_2632, signal_1014}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1004 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_2649, signal_2648, signal_2647, signal_1019}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1005 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_2652, signal_2651, signal_2650, signal_1020}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1006 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_2655, signal_2654, signal_2653, signal_1021}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1007 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_2658, signal_2657, signal_2656, signal_1022}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1008 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2469, signal_2468, signal_2467, signal_959}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_2661, signal_2660, signal_2659, signal_1023}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1009 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_2664, signal_2663, signal_2662, signal_1024}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1010 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_2667, signal_2666, signal_2665, signal_1025}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1011 ( .a ({signal_2457, signal_2456, signal_2455, signal_955}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_2670, signal_2669, signal_2668, signal_1026}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1012 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_2673, signal_2672, signal_2671, signal_1027}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1013 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_2676, signal_2675, signal_2674, signal_1028}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1014 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_2679, signal_2678, signal_2677, signal_1029}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1015 ( .a ({signal_2460, signal_2459, signal_2458, signal_956}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_2682, signal_2681, signal_2680, signal_1030}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1033 ( .a ({signal_2601, signal_2600, signal_2599, signal_1003}), .b ({signal_2736, signal_2735, signal_2734, signal_1048}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1040 ( .a ({signal_2634, signal_2633, signal_2632, signal_1014}), .b ({signal_2757, signal_2756, signal_2755, signal_1055}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1044 ( .a ({signal_2652, signal_2651, signal_2650, signal_1020}), .b ({signal_2769, signal_2768, signal_2767, signal_1059}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1045 ( .a ({signal_2661, signal_2660, signal_2659, signal_1023}), .b ({signal_2772, signal_2771, signal_2770, signal_1060}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1046 ( .a ({signal_2667, signal_2666, signal_2665, signal_1025}), .b ({signal_2775, signal_2774, signal_2773, signal_1061}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1047 ( .a ({signal_2670, signal_2669, signal_2668, signal_1026}), .b ({signal_2778, signal_2777, signal_2776, signal_1062}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1048 ( .a ({signal_2673, signal_2672, signal_2671, signal_1027}), .b ({signal_2781, signal_2780, signal_2779, signal_1063}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1049 ( .a ({signal_2676, signal_2675, signal_2674, signal_1028}), .b ({signal_2784, signal_2783, signal_2782, signal_1064}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1050 ( .a ({signal_2679, signal_2678, signal_2677, signal_1029}), .b ({signal_2787, signal_2786, signal_2785, signal_1065}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1051 ( .a ({signal_2682, signal_2681, signal_2680, signal_1030}), .b ({signal_2790, signal_2789, signal_2788, signal_1066}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1052 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2529, signal_2528, signal_2527, signal_979}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_2793, signal_2792, signal_2791, signal_1067}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1053 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_2796, signal_2795, signal_2794, signal_1068}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1054 ( .a ({signal_2493, signal_2492, signal_2491, signal_967}), .b ({signal_2496, signal_2495, signal_2494, signal_968}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_2799, signal_2798, signal_2797, signal_1069}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1055 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2490, signal_2489, signal_2488, signal_966}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_2802, signal_2801, signal_2800, signal_1070}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1056 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_2805, signal_2804, signal_2803, signal_1071}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1057 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_2808, signal_2807, signal_2806, signal_1072}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1058 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_2811, signal_2810, signal_2809, signal_1073}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1059 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2535, signal_2534, signal_2533, signal_981}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_2814, signal_2813, signal_2812, signal_1074}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1060 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_2817, signal_2816, signal_2815, signal_1075}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1061 ( .a ({signal_2574, signal_2573, signal_2572, signal_994}), .b ({signal_2589, signal_2588, signal_2587, signal_999}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_2820, signal_2819, signal_2818, signal_1076}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1062 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2529, signal_2528, signal_2527, signal_979}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_2823, signal_2822, signal_2821, signal_1077}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1063 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_2826, signal_2825, signal_2824, signal_1078}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1064 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2598, signal_2597, signal_2596, signal_1002}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_2829, signal_2828, signal_2827, signal_1079}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1065 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_2832, signal_2831, signal_2830, signal_1080}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1066 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_2835, signal_2834, signal_2833, signal_1081}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1067 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2547, signal_2546, signal_2545, signal_985}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_2838, signal_2837, signal_2836, signal_1082}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1068 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_2841, signal_2840, signal_2839, signal_1083}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1069 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_2844, signal_2843, signal_2842, signal_1084}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1070 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2586, signal_2585, signal_2584, signal_998}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_2847, signal_2846, signal_2845, signal_1085}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1071 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_2850, signal_2849, signal_2848, signal_1086}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1072 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_2853, signal_2852, signal_2851, signal_1087}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1073 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2544, signal_2543, signal_2542, signal_984}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_2856, signal_2855, signal_2854, signal_1088}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1074 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_2859, signal_2858, signal_2857, signal_1089}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1075 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_2862, signal_2861, signal_2860, signal_1090}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1076 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_2865, signal_2864, signal_2863, signal_1091}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1077 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_2868, signal_2867, signal_2866, signal_1092}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1078 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_2871, signal_2870, signal_2869, signal_1093}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1079 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_2874, signal_2873, signal_2872, signal_1094}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1080 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_2877, signal_2876, signal_2875, signal_1095}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1081 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_2880, signal_2879, signal_2878, signal_1096}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1082 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_2883, signal_2882, signal_2881, signal_1097}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1083 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2535, signal_2534, signal_2533, signal_981}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_2886, signal_2885, signal_2884, signal_1098}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1084 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_2889, signal_2888, signal_2887, signal_1099}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1086 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_2895, signal_2894, signal_2893, signal_1101}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1087 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2538, signal_2537, signal_2536, signal_982}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_2898, signal_2897, signal_2896, signal_1102}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1088 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_2901, signal_2900, signal_2899, signal_1103}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1089 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_2904, signal_2903, signal_2902, signal_1104}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1090 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_2907, signal_2906, signal_2905, signal_1105}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1091 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2640, signal_2639, signal_2638, signal_1016}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_2910, signal_2909, signal_2908, signal_1106}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1092 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_2913, signal_2912, signal_2911, signal_1107}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1093 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_2916, signal_2915, signal_2914, signal_1108}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1094 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_2919, signal_2918, signal_2917, signal_1109}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1095 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_2922, signal_2921, signal_2920, signal_1110}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1096 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_2925, signal_2924, signal_2923, signal_1111}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1097 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2631, signal_2630, signal_2629, signal_1013}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_2928, signal_2927, signal_2926, signal_1112}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1098 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_2931, signal_2930, signal_2929, signal_1113}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1099 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_2934, signal_2933, signal_2932, signal_1114}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1100 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_2937, signal_2936, signal_2935, signal_1115}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1101 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_2940, signal_2939, signal_2938, signal_1116}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1102 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_2943, signal_2942, signal_2941, signal_1117}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1103 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2598, signal_2597, signal_2596, signal_1002}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_2946, signal_2945, signal_2944, signal_1118}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1104 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_2949, signal_2948, signal_2947, signal_1119}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1105 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_2952, signal_2951, signal_2950, signal_1120}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1106 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_2955, signal_2954, signal_2953, signal_1121}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1107 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2646, signal_2645, signal_2644, signal_1018}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_2958, signal_2957, signal_2956, signal_1122}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1108 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_2961, signal_2960, signal_2959, signal_1123}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1109 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2589, signal_2588, signal_2587, signal_999}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_2964, signal_2963, signal_2962, signal_1124}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1110 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_2967, signal_2966, signal_2965, signal_1125}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1111 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_2970, signal_2969, signal_2968, signal_1126}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1112 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2460, signal_2459, signal_2458, signal_956}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_2973, signal_2972, signal_2971, signal_1127}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1113 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2481, signal_2480, signal_2479, signal_963}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_2976, signal_2975, signal_2974, signal_1128}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1114 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2640, signal_2639, signal_2638, signal_1016}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_2979, signal_2978, signal_2977, signal_1129}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1115 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_2982, signal_2981, signal_2980, signal_1130}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1116 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_2985, signal_2984, signal_2983, signal_1131}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1117 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2550, signal_2549, signal_2548, signal_986}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_2988, signal_2987, signal_2986, signal_1132}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1118 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2562, signal_2561, signal_2560, signal_990}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_2991, signal_2990, signal_2989, signal_1133}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1119 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_2994, signal_2993, signal_2992, signal_1134}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1120 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_2997, signal_2996, signal_2995, signal_1135}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1121 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_3000, signal_2999, signal_2998, signal_1136}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1122 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2577, signal_2576, signal_2575, signal_995}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_3003, signal_3002, signal_3001, signal_1137}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1123 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_3006, signal_3005, signal_3004, signal_1138}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1125 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_3012, signal_3011, signal_3010, signal_1140}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1126 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_3015, signal_3014, signal_3013, signal_1141}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1127 ( .a ({signal_2466, signal_2465, signal_2464, signal_958}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_3018, signal_3017, signal_3016, signal_1142}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1128 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_3021, signal_3020, signal_3019, signal_1143}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1129 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_3024, signal_3023, signal_3022, signal_1144}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1130 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_3027, signal_3026, signal_3025, signal_1145}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1131 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2610, signal_2609, signal_2608, signal_1006}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_3030, signal_3029, signal_3028, signal_1146}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1133 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_3036, signal_3035, signal_3034, signal_1148}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1134 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_3039, signal_3038, signal_3037, signal_1149}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1135 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_3042, signal_3041, signal_3040, signal_1150}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1136 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_3045, signal_3044, signal_3043, signal_1151}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1137 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_3048, signal_3047, signal_3046, signal_1152}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1138 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_3051, signal_3050, signal_3049, signal_1153}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1139 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_3054, signal_3053, signal_3052, signal_1154}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1141 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_3060, signal_3059, signal_3058, signal_1156}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1142 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_3063, signal_3062, signal_3061, signal_1157}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1143 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_3066, signal_3065, signal_3064, signal_1158}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1144 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2463, signal_2462, signal_2461, signal_957}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_3069, signal_3068, signal_3067, signal_1159}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1145 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_3072, signal_3071, signal_3070, signal_1160}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1146 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_3075, signal_3074, signal_3073, signal_1161}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1147 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_3078, signal_3077, signal_3076, signal_1162}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1148 ( .a ({signal_2490, signal_2489, signal_2488, signal_966}), .b ({signal_2511, signal_2510, signal_2509, signal_973}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_3081, signal_3080, signal_3079, signal_1163}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1149 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_3084, signal_3083, signal_3082, signal_1164}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1150 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2625, signal_2624, signal_2623, signal_1011}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_3087, signal_3086, signal_3085, signal_1165}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1151 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_3090, signal_3089, signal_3088, signal_1166}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1152 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_3093, signal_3092, signal_3091, signal_1167}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1153 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_3096, signal_3095, signal_3094, signal_1168}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1154 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_3099, signal_3098, signal_3097, signal_1169}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1156 ( .a ({signal_2610, signal_2609, signal_2608, signal_1006}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_3105, signal_3104, signal_3103, signal_1171}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1157 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_3108, signal_3107, signal_3106, signal_1172}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1158 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_3111, signal_3110, signal_3109, signal_1173}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1159 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_3114, signal_3113, signal_3112, signal_1174}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1160 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_3117, signal_3116, signal_3115, signal_1175}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1161 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_3120, signal_3119, signal_3118, signal_1176}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1162 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_3123, signal_3122, signal_3121, signal_1177}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1163 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_3126, signal_3125, signal_3124, signal_1178}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1164 ( .a ({signal_2490, signal_2489, signal_2488, signal_966}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_3129, signal_3128, signal_3127, signal_1179}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1165 ( .a ({signal_2505, signal_2504, signal_2503, signal_971}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_3132, signal_3131, signal_3130, signal_1180}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1166 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_3135, signal_3134, signal_3133, signal_1181}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1167 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_3138, signal_3137, signal_3136, signal_1182}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1168 ( .a ({signal_2457, signal_2456, signal_2455, signal_955}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_3141, signal_3140, signal_3139, signal_1183}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1169 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_3144, signal_3143, signal_3142, signal_1184}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1170 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_3147, signal_3146, signal_3145, signal_1185}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1171 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_3150, signal_3149, signal_3148, signal_1186}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1172 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2577, signal_2576, signal_2575, signal_995}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_3153, signal_3152, signal_3151, signal_1187}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1174 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2544, signal_2543, signal_2542, signal_984}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_3159, signal_3158, signal_3157, signal_1189}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1175 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_3162, signal_3161, signal_3160, signal_1190}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1176 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_3165, signal_3164, signal_3163, signal_1191}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1177 ( .a ({signal_2580, signal_2579, signal_2578, signal_996}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_3168, signal_3167, signal_3166, signal_1192}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1178 ( .a ({signal_2499, signal_2498, signal_2497, signal_969}), .b ({signal_2520, signal_2519, signal_2518, signal_976}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_3171, signal_3170, signal_3169, signal_1193}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1179 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_3174, signal_3173, signal_3172, signal_1194}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1180 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_2463, signal_2462, signal_2461, signal_957}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_3177, signal_3176, signal_3175, signal_1195}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1181 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_3180, signal_3179, signal_3178, signal_1196}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1182 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_3183, signal_3182, signal_3181, signal_1197}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1183 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_3186, signal_3185, signal_3184, signal_1198}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1185 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_3192, signal_3191, signal_3190, signal_1200}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1186 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_3195, signal_3194, signal_3193, signal_1201}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1187 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2547, signal_2546, signal_2545, signal_985}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_3198, signal_3197, signal_3196, signal_1202}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1188 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2469, signal_2468, signal_2467, signal_959}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_3201, signal_3200, signal_3199, signal_1203}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1191 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2553, signal_2552, signal_2551, signal_987}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_3210, signal_3209, signal_3208, signal_1206}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1192 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_3213, signal_3212, signal_3211, signal_1207}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1193 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_3216, signal_3215, signal_3214, signal_1208}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1194 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_3219, signal_3218, signal_3217, signal_1209}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1195 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_3222, signal_3221, signal_3220, signal_1210}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1196 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_3225, signal_3224, signal_3223, signal_1211}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1197 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2550, signal_2549, signal_2548, signal_986}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_3228, signal_3227, signal_3226, signal_1212}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1199 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_3234, signal_3233, signal_3232, signal_1214}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1200 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_3237, signal_3236, signal_3235, signal_1215}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1201 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2586, signal_2585, signal_2584, signal_998}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_3240, signal_3239, signal_3238, signal_1216}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1202 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({signal_3243, signal_3242, signal_3241, signal_1217}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1203 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({signal_3246, signal_3245, signal_3244, signal_1218}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1204 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({signal_3249, signal_3248, signal_3247, signal_1219}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1205 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({signal_3252, signal_3251, signal_3250, signal_1220}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1206 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_3255, signal_3254, signal_3253, signal_1221}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1208 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({signal_3261, signal_3260, signal_3259, signal_1223}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1210 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2502, signal_2501, signal_2500, signal_970}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({signal_3267, signal_3266, signal_3265, signal_1225}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1213 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2526, signal_2525, signal_2524, signal_978}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({signal_3276, signal_3275, signal_3274, signal_1228}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1214 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({signal_3279, signal_3278, signal_3277, signal_1229}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1215 ( .a ({signal_2799, signal_2798, signal_2797, signal_1069}), .b ({signal_3282, signal_3281, signal_3280, signal_1230}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1216 ( .a ({signal_2802, signal_2801, signal_2800, signal_1070}), .b ({signal_3285, signal_3284, signal_3283, signal_1231}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1217 ( .a ({signal_2808, signal_2807, signal_2806, signal_1072}), .b ({signal_3288, signal_3287, signal_3286, signal_1232}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1218 ( .a ({signal_2811, signal_2810, signal_2809, signal_1073}), .b ({signal_3291, signal_3290, signal_3289, signal_1233}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1219 ( .a ({signal_2814, signal_2813, signal_2812, signal_1074}), .b ({signal_3294, signal_3293, signal_3292, signal_1234}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1220 ( .a ({signal_2817, signal_2816, signal_2815, signal_1075}), .b ({signal_3297, signal_3296, signal_3295, signal_1235}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1221 ( .a ({signal_2820, signal_2819, signal_2818, signal_1076}), .b ({signal_3300, signal_3299, signal_3298, signal_1236}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1222 ( .a ({signal_2823, signal_2822, signal_2821, signal_1077}), .b ({signal_3303, signal_3302, signal_3301, signal_1237}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1223 ( .a ({signal_2826, signal_2825, signal_2824, signal_1078}), .b ({signal_3306, signal_3305, signal_3304, signal_1238}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1224 ( .a ({signal_2829, signal_2828, signal_2827, signal_1079}), .b ({signal_3309, signal_3308, signal_3307, signal_1239}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1225 ( .a ({signal_2832, signal_2831, signal_2830, signal_1080}), .b ({signal_3312, signal_3311, signal_3310, signal_1240}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1226 ( .a ({signal_2835, signal_2834, signal_2833, signal_1081}), .b ({signal_3315, signal_3314, signal_3313, signal_1241}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1227 ( .a ({signal_2838, signal_2837, signal_2836, signal_1082}), .b ({signal_3318, signal_3317, signal_3316, signal_1242}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1228 ( .a ({signal_2841, signal_2840, signal_2839, signal_1083}), .b ({signal_3321, signal_3320, signal_3319, signal_1243}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1229 ( .a ({signal_2844, signal_2843, signal_2842, signal_1084}), .b ({signal_3324, signal_3323, signal_3322, signal_1244}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1230 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_3327, signal_3326, signal_3325, signal_1245}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1231 ( .a ({signal_2853, signal_2852, signal_2851, signal_1087}), .b ({signal_3330, signal_3329, signal_3328, signal_1246}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1232 ( .a ({signal_2856, signal_2855, signal_2854, signal_1088}), .b ({signal_3333, signal_3332, signal_3331, signal_1247}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1233 ( .a ({signal_2862, signal_2861, signal_2860, signal_1090}), .b ({signal_3336, signal_3335, signal_3334, signal_1248}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1234 ( .a ({signal_2865, signal_2864, signal_2863, signal_1091}), .b ({signal_3339, signal_3338, signal_3337, signal_1249}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1235 ( .a ({signal_2868, signal_2867, signal_2866, signal_1092}), .b ({signal_3342, signal_3341, signal_3340, signal_1250}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1236 ( .a ({signal_2871, signal_2870, signal_2869, signal_1093}), .b ({signal_3345, signal_3344, signal_3343, signal_1251}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1237 ( .a ({signal_2874, signal_2873, signal_2872, signal_1094}), .b ({signal_3348, signal_3347, signal_3346, signal_1252}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1238 ( .a ({signal_2877, signal_2876, signal_2875, signal_1095}), .b ({signal_3351, signal_3350, signal_3349, signal_1253}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1239 ( .a ({signal_2880, signal_2879, signal_2878, signal_1096}), .b ({signal_3354, signal_3353, signal_3352, signal_1254}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1240 ( .a ({signal_2883, signal_2882, signal_2881, signal_1097}), .b ({signal_3357, signal_3356, signal_3355, signal_1255}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1241 ( .a ({signal_2886, signal_2885, signal_2884, signal_1098}), .b ({signal_3360, signal_3359, signal_3358, signal_1256}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1242 ( .a ({signal_2889, signal_2888, signal_2887, signal_1099}), .b ({signal_3363, signal_3362, signal_3361, signal_1257}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1244 ( .a ({signal_2895, signal_2894, signal_2893, signal_1101}), .b ({signal_3369, signal_3368, signal_3367, signal_1259}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1245 ( .a ({signal_2901, signal_2900, signal_2899, signal_1103}), .b ({signal_3372, signal_3371, signal_3370, signal_1260}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1246 ( .a ({signal_2907, signal_2906, signal_2905, signal_1105}), .b ({signal_3375, signal_3374, signal_3373, signal_1261}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1247 ( .a ({signal_2910, signal_2909, signal_2908, signal_1106}), .b ({signal_3378, signal_3377, signal_3376, signal_1262}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1248 ( .a ({signal_2916, signal_2915, signal_2914, signal_1108}), .b ({signal_3381, signal_3380, signal_3379, signal_1263}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1249 ( .a ({signal_2919, signal_2918, signal_2917, signal_1109}), .b ({signal_3384, signal_3383, signal_3382, signal_1264}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1250 ( .a ({signal_2922, signal_2921, signal_2920, signal_1110}), .b ({signal_3387, signal_3386, signal_3385, signal_1265}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1251 ( .a ({signal_2925, signal_2924, signal_2923, signal_1111}), .b ({signal_3390, signal_3389, signal_3388, signal_1266}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1252 ( .a ({signal_2928, signal_2927, signal_2926, signal_1112}), .b ({signal_3393, signal_3392, signal_3391, signal_1267}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1253 ( .a ({signal_2931, signal_2930, signal_2929, signal_1113}), .b ({signal_3396, signal_3395, signal_3394, signal_1268}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1254 ( .a ({signal_2937, signal_2936, signal_2935, signal_1115}), .b ({signal_3399, signal_3398, signal_3397, signal_1269}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1255 ( .a ({signal_2940, signal_2939, signal_2938, signal_1116}), .b ({signal_3402, signal_3401, signal_3400, signal_1270}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1256 ( .a ({signal_2943, signal_2942, signal_2941, signal_1117}), .b ({signal_3405, signal_3404, signal_3403, signal_1271}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1257 ( .a ({signal_2946, signal_2945, signal_2944, signal_1118}), .b ({signal_3408, signal_3407, signal_3406, signal_1272}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1258 ( .a ({signal_2952, signal_2951, signal_2950, signal_1120}), .b ({signal_3411, signal_3410, signal_3409, signal_1273}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1259 ( .a ({signal_2955, signal_2954, signal_2953, signal_1121}), .b ({signal_3414, signal_3413, signal_3412, signal_1274}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1260 ( .a ({signal_2958, signal_2957, signal_2956, signal_1122}), .b ({signal_3417, signal_3416, signal_3415, signal_1275}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1261 ( .a ({signal_2964, signal_2963, signal_2962, signal_1124}), .b ({signal_3420, signal_3419, signal_3418, signal_1276}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1262 ( .a ({signal_2967, signal_2966, signal_2965, signal_1125}), .b ({signal_3423, signal_3422, signal_3421, signal_1277}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1263 ( .a ({signal_2970, signal_2969, signal_2968, signal_1126}), .b ({signal_3426, signal_3425, signal_3424, signal_1278}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1264 ( .a ({signal_2973, signal_2972, signal_2971, signal_1127}), .b ({signal_3429, signal_3428, signal_3427, signal_1279}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1265 ( .a ({signal_2979, signal_2978, signal_2977, signal_1129}), .b ({signal_3432, signal_3431, signal_3430, signal_1280}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1266 ( .a ({signal_2982, signal_2981, signal_2980, signal_1130}), .b ({signal_3435, signal_3434, signal_3433, signal_1281}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1267 ( .a ({signal_2985, signal_2984, signal_2983, signal_1131}), .b ({signal_3438, signal_3437, signal_3436, signal_1282}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1268 ( .a ({signal_2994, signal_2993, signal_2992, signal_1134}), .b ({signal_3441, signal_3440, signal_3439, signal_1283}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1269 ( .a ({signal_2997, signal_2996, signal_2995, signal_1135}), .b ({signal_3444, signal_3443, signal_3442, signal_1284}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1270 ( .a ({signal_3000, signal_2999, signal_2998, signal_1136}), .b ({signal_3447, signal_3446, signal_3445, signal_1285}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1271 ( .a ({signal_3003, signal_3002, signal_3001, signal_1137}), .b ({signal_3450, signal_3449, signal_3448, signal_1286}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1273 ( .a ({signal_3015, signal_3014, signal_3013, signal_1141}), .b ({signal_3456, signal_3455, signal_3454, signal_1288}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1274 ( .a ({signal_3021, signal_3020, signal_3019, signal_1143}), .b ({signal_3459, signal_3458, signal_3457, signal_1289}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1275 ( .a ({signal_3024, signal_3023, signal_3022, signal_1144}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1276 ( .a ({signal_3030, signal_3029, signal_3028, signal_1146}), .b ({signal_3465, signal_3464, signal_3463, signal_1291}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1278 ( .a ({signal_3036, signal_3035, signal_3034, signal_1148}), .b ({signal_3471, signal_3470, signal_3469, signal_1293}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1279 ( .a ({signal_3039, signal_3038, signal_3037, signal_1149}), .b ({signal_3474, signal_3473, signal_3472, signal_1294}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1280 ( .a ({signal_3042, signal_3041, signal_3040, signal_1150}), .b ({signal_3477, signal_3476, signal_3475, signal_1295}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1281 ( .a ({signal_3048, signal_3047, signal_3046, signal_1152}), .b ({signal_3480, signal_3479, signal_3478, signal_1296}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1282 ( .a ({signal_3051, signal_3050, signal_3049, signal_1153}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1283 ( .a ({signal_3054, signal_3053, signal_3052, signal_1154}), .b ({signal_3486, signal_3485, signal_3484, signal_1298}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1285 ( .a ({signal_3060, signal_3059, signal_3058, signal_1156}), .b ({signal_3492, signal_3491, signal_3490, signal_1300}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1286 ( .a ({signal_3063, signal_3062, signal_3061, signal_1157}), .b ({signal_3495, signal_3494, signal_3493, signal_1301}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1287 ( .a ({signal_3069, signal_3068, signal_3067, signal_1159}), .b ({signal_3498, signal_3497, signal_3496, signal_1302}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1288 ( .a ({signal_3072, signal_3071, signal_3070, signal_1160}), .b ({signal_3501, signal_3500, signal_3499, signal_1303}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1289 ( .a ({signal_3075, signal_3074, signal_3073, signal_1161}), .b ({signal_3504, signal_3503, signal_3502, signal_1304}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1290 ( .a ({signal_3078, signal_3077, signal_3076, signal_1162}), .b ({signal_3507, signal_3506, signal_3505, signal_1305}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1291 ( .a ({signal_3081, signal_3080, signal_3079, signal_1163}), .b ({signal_3510, signal_3509, signal_3508, signal_1306}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1292 ( .a ({signal_3084, signal_3083, signal_3082, signal_1164}), .b ({signal_3513, signal_3512, signal_3511, signal_1307}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1293 ( .a ({signal_3087, signal_3086, signal_3085, signal_1165}), .b ({signal_3516, signal_3515, signal_3514, signal_1308}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1294 ( .a ({signal_3090, signal_3089, signal_3088, signal_1166}), .b ({signal_3519, signal_3518, signal_3517, signal_1309}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1295 ( .a ({signal_3093, signal_3092, signal_3091, signal_1167}), .b ({signal_3522, signal_3521, signal_3520, signal_1310}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1296 ( .a ({signal_3099, signal_3098, signal_3097, signal_1169}), .b ({signal_3525, signal_3524, signal_3523, signal_1311}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1298 ( .a ({signal_3105, signal_3104, signal_3103, signal_1171}), .b ({signal_3531, signal_3530, signal_3529, signal_1313}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1299 ( .a ({signal_3108, signal_3107, signal_3106, signal_1172}), .b ({signal_3534, signal_3533, signal_3532, signal_1314}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1300 ( .a ({signal_3111, signal_3110, signal_3109, signal_1173}), .b ({signal_3537, signal_3536, signal_3535, signal_1315}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1301 ( .a ({signal_3114, signal_3113, signal_3112, signal_1174}), .b ({signal_3540, signal_3539, signal_3538, signal_1316}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1302 ( .a ({signal_3117, signal_3116, signal_3115, signal_1175}), .b ({signal_3543, signal_3542, signal_3541, signal_1317}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1303 ( .a ({signal_3120, signal_3119, signal_3118, signal_1176}), .b ({signal_3546, signal_3545, signal_3544, signal_1318}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1304 ( .a ({signal_3123, signal_3122, signal_3121, signal_1177}), .b ({signal_3549, signal_3548, signal_3547, signal_1319}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1305 ( .a ({signal_3129, signal_3128, signal_3127, signal_1179}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1306 ( .a ({signal_3132, signal_3131, signal_3130, signal_1180}), .b ({signal_3555, signal_3554, signal_3553, signal_1321}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1307 ( .a ({signal_3135, signal_3134, signal_3133, signal_1181}), .b ({signal_3558, signal_3557, signal_3556, signal_1322}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1308 ( .a ({signal_3138, signal_3137, signal_3136, signal_1182}), .b ({signal_3561, signal_3560, signal_3559, signal_1323}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1309 ( .a ({signal_3141, signal_3140, signal_3139, signal_1183}), .b ({signal_3564, signal_3563, signal_3562, signal_1324}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1310 ( .a ({signal_3144, signal_3143, signal_3142, signal_1184}), .b ({signal_3567, signal_3566, signal_3565, signal_1325}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1311 ( .a ({signal_3147, signal_3146, signal_3145, signal_1185}), .b ({signal_3570, signal_3569, signal_3568, signal_1326}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1312 ( .a ({signal_3150, signal_3149, signal_3148, signal_1186}), .b ({signal_3573, signal_3572, signal_3571, signal_1327}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1313 ( .a ({signal_3153, signal_3152, signal_3151, signal_1187}), .b ({signal_3576, signal_3575, signal_3574, signal_1328}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1315 ( .a ({signal_3159, signal_3158, signal_3157, signal_1189}), .b ({signal_3582, signal_3581, signal_3580, signal_1330}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1316 ( .a ({signal_3165, signal_3164, signal_3163, signal_1191}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1317 ( .a ({signal_3168, signal_3167, signal_3166, signal_1192}), .b ({signal_3588, signal_3587, signal_3586, signal_1332}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1318 ( .a ({signal_3171, signal_3170, signal_3169, signal_1193}), .b ({signal_3591, signal_3590, signal_3589, signal_1333}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1319 ( .a ({signal_3174, signal_3173, signal_3172, signal_1194}), .b ({signal_3594, signal_3593, signal_3592, signal_1334}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1320 ( .a ({signal_3177, signal_3176, signal_3175, signal_1195}), .b ({signal_3597, signal_3596, signal_3595, signal_1335}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1321 ( .a ({signal_3180, signal_3179, signal_3178, signal_1196}), .b ({signal_3600, signal_3599, signal_3598, signal_1336}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1322 ( .a ({signal_3183, signal_3182, signal_3181, signal_1197}), .b ({signal_3603, signal_3602, signal_3601, signal_1337}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1324 ( .a ({signal_3192, signal_3191, signal_3190, signal_1200}), .b ({signal_3609, signal_3608, signal_3607, signal_1339}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1325 ( .a ({signal_3195, signal_3194, signal_3193, signal_1201}), .b ({signal_3612, signal_3611, signal_3610, signal_1340}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1326 ( .a ({signal_3198, signal_3197, signal_3196, signal_1202}), .b ({signal_3615, signal_3614, signal_3613, signal_1341}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1327 ( .a ({signal_3201, signal_3200, signal_3199, signal_1203}), .b ({signal_3618, signal_3617, signal_3616, signal_1342}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1330 ( .a ({signal_3213, signal_3212, signal_3211, signal_1207}), .b ({signal_3627, signal_3626, signal_3625, signal_1345}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1331 ( .a ({signal_3219, signal_3218, signal_3217, signal_1209}), .b ({signal_3630, signal_3629, signal_3628, signal_1346}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1332 ( .a ({signal_3222, signal_3221, signal_3220, signal_1210}), .b ({signal_3633, signal_3632, signal_3631, signal_1347}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1333 ( .a ({signal_3225, signal_3224, signal_3223, signal_1211}), .b ({signal_3636, signal_3635, signal_3634, signal_1348}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1334 ( .a ({signal_3228, signal_3227, signal_3226, signal_1212}), .b ({signal_3639, signal_3638, signal_3637, signal_1349}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1336 ( .a ({signal_3234, signal_3233, signal_3232, signal_1214}), .b ({signal_3645, signal_3644, signal_3643, signal_1351}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1337 ( .a ({signal_3237, signal_3236, signal_3235, signal_1215}), .b ({signal_3648, signal_3647, signal_3646, signal_1352}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1338 ( .a ({signal_3240, signal_3239, signal_3238, signal_1216}), .b ({signal_3651, signal_3650, signal_3649, signal_1353}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1339 ( .a ({signal_3246, signal_3245, signal_3244, signal_1218}), .b ({signal_3654, signal_3653, signal_3652, signal_1354}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1340 ( .a ({signal_3249, signal_3248, signal_3247, signal_1219}), .b ({signal_3657, signal_3656, signal_3655, signal_1355}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1341 ( .a ({signal_3252, signal_3251, signal_3250, signal_1220}), .b ({signal_3660, signal_3659, signal_3658, signal_1356}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1342 ( .a ({signal_3255, signal_3254, signal_3253, signal_1221}), .b ({signal_3663, signal_3662, signal_3661, signal_1357}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1344 ( .a ({signal_3261, signal_3260, signal_3259, signal_1223}), .b ({signal_3669, signal_3668, signal_3667, signal_1359}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1346 ( .a ({signal_3267, signal_3266, signal_3265, signal_1225}), .b ({signal_3675, signal_3674, signal_3673, signal_1361}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1349 ( .a ({signal_3276, signal_3275, signal_3274, signal_1228}), .b ({signal_3684, signal_3683, signal_3682, signal_1364}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1350 ( .a ({signal_3279, signal_3278, signal_3277, signal_1229}), .b ({signal_3687, signal_3686, signal_3685, signal_1365}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1353 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_3696, signal_3695, signal_3694, signal_1368}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1354 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2718, signal_2717, signal_2716, signal_1042}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({signal_3699, signal_3698, signal_3697, signal_1369}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1355 ( .a ({signal_2685, signal_2684, signal_2683, signal_1031}), .b ({signal_2766, signal_2765, signal_2764, signal_1058}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({signal_3702, signal_3701, signal_3700, signal_1370}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1356 ( .a ({signal_2727, signal_2726, signal_2725, signal_1045}), .b ({signal_2763, signal_2762, signal_2761, signal_1057}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({signal_3705, signal_3704, signal_3703, signal_1371}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1357 ( .a ({signal_2700, signal_2699, signal_2698, signal_1036}), .b ({signal_2703, signal_2702, signal_2701, signal_1037}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({signal_3708, signal_3707, signal_3706, signal_1372}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1360 ( .a ({signal_2700, signal_2699, signal_2698, signal_1036}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_3717, signal_3716, signal_3715, signal_1375}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1361 ( .a ({signal_2715, signal_2714, signal_2713, signal_1041}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({signal_3720, signal_3719, signal_3718, signal_1376}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1362 ( .a ({signal_2745, signal_2744, signal_2743, signal_1051}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({signal_3723, signal_3722, signal_3721, signal_1377}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1365 ( .a ({signal_2685, signal_2684, signal_2683, signal_1031}), .b ({signal_2724, signal_2723, signal_2722, signal_1044}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({signal_3732, signal_3731, signal_3730, signal_1380}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1366 ( .a ({signal_2688, signal_2687, signal_2686, signal_1032}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({signal_3735, signal_3734, signal_3733, signal_1381}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1367 ( .a ({signal_2718, signal_2717, signal_2716, signal_1042}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_3738, signal_3737, signal_3736, signal_1382}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1368 ( .a ({signal_2703, signal_2702, signal_2701, signal_1037}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({signal_3741, signal_3740, signal_3739, signal_1383}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1369 ( .a ({signal_2514, signal_2513, signal_2512, signal_974}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({signal_3744, signal_3743, signal_3742, signal_1384}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1375 ( .a ({signal_2712, signal_2711, signal_2710, signal_1040}), .b ({signal_2760, signal_2759, signal_2758, signal_1056}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({signal_3762, signal_3761, signal_3760, signal_1390}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1376 ( .a ({signal_2727, signal_2726, signal_2725, signal_1045}), .b ({signal_2742, signal_2741, signal_2740, signal_1050}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({signal_3765, signal_3764, signal_3763, signal_1391}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1383 ( .a ({signal_2691, signal_2690, signal_2689, signal_1033}), .b ({signal_2697, signal_2696, signal_2695, signal_1035}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_3786, signal_3785, signal_3784, signal_1398}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1395 ( .a ({signal_2505, signal_2504, signal_2503, signal_971}), .b ({signal_2739, signal_2738, signal_2737, signal_1049}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({signal_3822, signal_3821, signal_3820, signal_1410}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1396 ( .a ({signal_2688, signal_2687, signal_2686, signal_1032}), .b ({signal_2733, signal_2732, signal_2731, signal_1047}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({signal_3825, signal_3824, signal_3823, signal_1411}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1401 ( .a ({signal_2493, signal_2492, signal_2491, signal_967}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({signal_3840, signal_3839, signal_3838, signal_1416}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1402 ( .a ({signal_2742, signal_2741, signal_2740, signal_1050}), .b ({signal_2517, signal_2516, signal_2515, signal_975}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({signal_3843, signal_3842, signal_3841, signal_1417}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1403 ( .a ({signal_2508, signal_2507, signal_2506, signal_972}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_3846, signal_3845, signal_3844, signal_1418}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1407 ( .a ({signal_2706, signal_2705, signal_2704, signal_1038}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({signal_3858, signal_3857, signal_3856, signal_1422}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1408 ( .a ({signal_2712, signal_2711, signal_2710, signal_1040}), .b ({signal_2517, signal_2516, signal_2515, signal_975}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({signal_3861, signal_3860, signal_3859, signal_1423}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1492 ( .a ({signal_3696, signal_3695, signal_3694, signal_1368}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1493 ( .a ({signal_3699, signal_3698, signal_3697, signal_1369}), .b ({signal_4116, signal_4115, signal_4114, signal_1508}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1494 ( .a ({signal_3702, signal_3701, signal_3700, signal_1370}), .b ({signal_4119, signal_4118, signal_4117, signal_1509}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1495 ( .a ({signal_3705, signal_3704, signal_3703, signal_1371}), .b ({signal_4122, signal_4121, signal_4120, signal_1510}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1496 ( .a ({signal_3708, signal_3707, signal_3706, signal_1372}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1499 ( .a ({signal_3717, signal_3716, signal_3715, signal_1375}), .b ({signal_4134, signal_4133, signal_4132, signal_1514}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1500 ( .a ({signal_3720, signal_3719, signal_3718, signal_1376}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1501 ( .a ({signal_3723, signal_3722, signal_3721, signal_1377}), .b ({signal_4140, signal_4139, signal_4138, signal_1516}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1504 ( .a ({signal_3732, signal_3731, signal_3730, signal_1380}), .b ({signal_4149, signal_4148, signal_4147, signal_1519}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1505 ( .a ({signal_3735, signal_3734, signal_3733, signal_1381}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1506 ( .a ({signal_3738, signal_3737, signal_3736, signal_1382}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1507 ( .a ({signal_3744, signal_3743, signal_3742, signal_1384}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1513 ( .a ({signal_3765, signal_3764, signal_3763, signal_1391}), .b ({signal_4176, signal_4175, signal_4174, signal_1528}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1520 ( .a ({signal_3786, signal_3785, signal_3784, signal_1398}), .b ({signal_4197, signal_4196, signal_4195, signal_1535}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1532 ( .a ({signal_3822, signal_3821, signal_3820, signal_1410}), .b ({signal_4233, signal_4232, signal_4231, signal_1547}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1533 ( .a ({signal_3825, signal_3824, signal_3823, signal_1411}), .b ({signal_4236, signal_4235, signal_4234, signal_1548}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1538 ( .a ({signal_3840, signal_3839, signal_3838, signal_1416}), .b ({signal_4251, signal_4250, signal_4249, signal_1553}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1539 ( .a ({signal_3843, signal_3842, signal_3841, signal_1417}), .b ({signal_4254, signal_4253, signal_4252, signal_1554}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1543 ( .a ({signal_3858, signal_3857, signal_3856, signal_1422}), .b ({signal_4266, signal_4265, signal_4264, signal_1558}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1544 ( .a ({signal_3861, signal_3860, signal_3859, signal_1423}), .b ({signal_4269, signal_4268, signal_4267, signal_1559}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1085 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2634, signal_2633, signal_2632, signal_1014}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({signal_2892, signal_2891, signal_2890, signal_1100}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1124 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2649, signal_2648, signal_2647, signal_1019}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({signal_3009, signal_3008, signal_3007, signal_1139}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1132 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_3033, signal_3032, signal_3031, signal_1147}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1140 ( .a ({signal_2622, signal_2621, signal_2620, signal_1010}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({signal_3057, signal_3056, signal_3055, signal_1155}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1155 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({signal_3102, signal_3101, signal_3100, signal_1170}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1173 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({signal_3156, signal_3155, signal_3154, signal_1188}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1184 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({signal_3189, signal_3188, signal_3187, signal_1199}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1189 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_3204, signal_3203, signal_3202, signal_1204}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1190 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({signal_3207, signal_3206, signal_3205, signal_1205}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1198 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({signal_3231, signal_3230, signal_3229, signal_1213}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1207 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({signal_3258, signal_3257, signal_3256, signal_1222}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1209 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2670, signal_2669, signal_2668, signal_1026}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({signal_3264, signal_3263, signal_3262, signal_1224}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1211 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_3270, signal_3269, signal_3268, signal_1226}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1212 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({signal_3273, signal_3272, signal_3271, signal_1227}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1243 ( .a ({signal_2892, signal_2891, signal_2890, signal_1100}), .b ({signal_3366, signal_3365, signal_3364, signal_1258}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1272 ( .a ({signal_3009, signal_3008, signal_3007, signal_1139}), .b ({signal_3453, signal_3452, signal_3451, signal_1287}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1277 ( .a ({signal_3033, signal_3032, signal_3031, signal_1147}), .b ({signal_3468, signal_3467, signal_3466, signal_1292}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1284 ( .a ({signal_3057, signal_3056, signal_3055, signal_1155}), .b ({signal_3489, signal_3488, signal_3487, signal_1299}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1297 ( .a ({signal_3102, signal_3101, signal_3100, signal_1170}), .b ({signal_3528, signal_3527, signal_3526, signal_1312}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1314 ( .a ({signal_3156, signal_3155, signal_3154, signal_1188}), .b ({signal_3579, signal_3578, signal_3577, signal_1329}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1323 ( .a ({signal_3189, signal_3188, signal_3187, signal_1199}), .b ({signal_3606, signal_3605, signal_3604, signal_1338}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1328 ( .a ({signal_3204, signal_3203, signal_3202, signal_1204}), .b ({signal_3621, signal_3620, signal_3619, signal_1343}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1329 ( .a ({signal_3207, signal_3206, signal_3205, signal_1205}), .b ({signal_3624, signal_3623, signal_3622, signal_1344}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1335 ( .a ({signal_3231, signal_3230, signal_3229, signal_1213}), .b ({signal_3642, signal_3641, signal_3640, signal_1350}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1343 ( .a ({signal_3258, signal_3257, signal_3256, signal_1222}), .b ({signal_3666, signal_3665, signal_3664, signal_1358}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1345 ( .a ({signal_3264, signal_3263, signal_3262, signal_1224}), .b ({signal_3672, signal_3671, signal_3670, signal_1360}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1347 ( .a ({signal_3270, signal_3269, signal_3268, signal_1226}), .b ({signal_3678, signal_3677, signal_3676, signal_1362}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1348 ( .a ({signal_3273, signal_3272, signal_3271, signal_1227}), .b ({signal_3681, signal_3680, signal_3679, signal_1363}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1351 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2793, signal_2792, signal_2791, signal_1067}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({signal_3690, signal_3689, signal_3688, signal_1366}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1352 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2796, signal_2795, signal_2794, signal_1068}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({signal_3693, signal_3692, signal_3691, signal_1367}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1358 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2832, signal_2831, signal_2830, signal_1080}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({signal_3711, signal_3710, signal_3709, signal_1373}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1359 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2847, signal_2846, signal_2845, signal_1085}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_3714, signal_3713, signal_3712, signal_1374}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1363 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2859, signal_2858, signal_2857, signal_1089}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({signal_3726, signal_3725, signal_3724, signal_1378}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1364 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({signal_3729, signal_3728, signal_3727, signal_1379}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1370 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({signal_3747, signal_3746, signal_3745, signal_1385}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1371 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({signal_3750, signal_3749, signal_3748, signal_1386}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1372 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_3753, signal_3752, signal_3751, signal_1387}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1373 ( .a ({signal_2811, signal_2810, signal_2809, signal_1073}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({signal_3756, signal_3755, signal_3754, signal_1388}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1374 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2883, signal_2882, signal_2881, signal_1097}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({signal_3759, signal_3758, signal_3757, signal_1389}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1377 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2904, signal_2903, signal_2902, signal_1104}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({signal_3768, signal_3767, signal_3766, signal_1392}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1378 ( .a ({signal_2688, signal_2687, signal_2686, signal_1032}), .b ({signal_2826, signal_2825, signal_2824, signal_1078}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({signal_3771, signal_3770, signal_3769, signal_1393}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1379 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_3774, signal_3773, signal_3772, signal_1394}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1380 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2859, signal_2858, signal_2857, signal_1089}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({signal_3777, signal_3776, signal_3775, signal_1395}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1381 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({signal_3780, signal_3779, signal_3778, signal_1396}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1382 ( .a ({signal_2640, signal_2639, signal_2638, signal_1016}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({signal_3783, signal_3782, signal_3781, signal_1397}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1384 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2913, signal_2912, signal_2911, signal_1107}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({signal_3789, signal_3788, signal_3787, signal_1399}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1385 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_2868, signal_2867, signal_2866, signal_1092}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_3792, signal_3791, signal_3790, signal_1400}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1386 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2832, signal_2831, signal_2830, signal_1080}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({signal_3795, signal_3794, signal_3793, signal_1401}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1387 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2850, signal_2849, signal_2848, signal_1086}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({signal_3798, signal_3797, signal_3796, signal_1402}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1388 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2934, signal_2933, signal_2932, signal_1114}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({signal_3801, signal_3800, signal_3799, signal_1403}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1389 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_2916, signal_2915, signal_2914, signal_1108}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({signal_3804, signal_3803, signal_3802, signal_1404}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1390 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_3807, signal_3806, signal_3805, signal_1405}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1391 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2883, signal_2882, signal_2881, signal_1097}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({signal_3810, signal_3809, signal_3808, signal_1406}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1392 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({signal_3813, signal_3812, signal_3811, signal_1407}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1393 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({signal_3816, signal_3815, signal_3814, signal_1408}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1394 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2934, signal_2933, signal_2932, signal_1114}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({signal_3819, signal_3818, signal_3817, signal_1409}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1397 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2898, signal_2897, signal_2896, signal_1102}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_3828, signal_3827, signal_3826, signal_1412}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1398 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2961, signal_2960, signal_2959, signal_1123}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({signal_3831, signal_3830, signal_3829, signal_1413}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1399 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({signal_3834, signal_3833, signal_3832, signal_1414}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1400 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({signal_3837, signal_3836, signal_3835, signal_1415}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1404 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2826, signal_2825, signal_2824, signal_1078}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({signal_3849, signal_3848, signal_3847, signal_1419}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1405 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2898, signal_2897, signal_2896, signal_1102}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_3852, signal_3851, signal_3850, signal_1420}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1406 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2937, signal_2936, signal_2935, signal_1115}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({signal_3855, signal_3854, signal_3853, signal_1421}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1409 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({signal_3864, signal_3863, signal_3862, signal_1424}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1410 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2913, signal_2912, signal_2911, signal_1107}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({signal_3867, signal_3866, signal_3865, signal_1425}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1411 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2850, signal_2849, signal_2848, signal_1086}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({signal_3870, signal_3869, signal_3868, signal_1426}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1412 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2976, signal_2975, signal_2974, signal_1128}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_3873, signal_3872, signal_3871, signal_1427}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1413 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2808, signal_2807, signal_2806, signal_1072}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({signal_3876, signal_3875, signal_3874, signal_1428}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1414 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2991, signal_2990, signal_2989, signal_1133}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({signal_3879, signal_3878, signal_3877, signal_1429}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1415 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({signal_3882, signal_3881, signal_3880, signal_1430}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1416 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({signal_3006, signal_3005, signal_3004, signal_1138}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({signal_3885, signal_3884, signal_3883, signal_1431}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1417 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_3888, signal_3887, signal_3886, signal_1432}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1418 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_3012, signal_3011, signal_3010, signal_1140}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({signal_3891, signal_3890, signal_3889, signal_1433}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1419 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({signal_3894, signal_3893, signal_3892, signal_1434}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1420 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_3018, signal_3017, signal_3016, signal_1142}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({signal_3897, signal_3896, signal_3895, signal_1435}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1421 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({signal_3900, signal_3899, signal_3898, signal_1436}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1422 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_3903, signal_3902, signal_3901, signal_1437}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1423 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_3045, signal_3044, signal_3043, signal_1151}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({signal_3906, signal_3905, signal_3904, signal_1438}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1424 ( .a ({signal_2613, signal_2612, signal_2611, signal_1007}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({signal_3909, signal_3908, signal_3907, signal_1439}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1425 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_3060, signal_3059, signal_3058, signal_1156}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({signal_3912, signal_3911, signal_3910, signal_1440}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1426 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({signal_3915, signal_3914, signal_3913, signal_1441}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1427 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_3918, signal_3917, signal_3916, signal_1442}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1428 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({signal_3921, signal_3920, signal_3919, signal_1443}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1429 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_3090, signal_3089, signal_3088, signal_1166}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({signal_3924, signal_3923, signal_3922, signal_1444}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1430 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({signal_3927, signal_3926, signal_3925, signal_1445}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1431 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_3096, signal_3095, signal_3094, signal_1168}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({signal_3930, signal_3929, signal_3928, signal_1446}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1432 ( .a ({signal_2658, signal_2657, signal_2656, signal_1022}), .b ({signal_3018, signal_3017, signal_3016, signal_1142}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_3933, signal_3932, signal_3931, signal_1447}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1433 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_3000, signal_2999, signal_2998, signal_1136}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({signal_3936, signal_3935, signal_3934, signal_1448}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1434 ( .a ({signal_3021, signal_3020, signal_3019, signal_1143}), .b ({signal_3027, signal_3026, signal_3025, signal_1145}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({signal_3939, signal_3938, signal_3937, signal_1449}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1435 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_3090, signal_3089, signal_3088, signal_1166}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({signal_3942, signal_3941, signal_3940, signal_1450}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1436 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({signal_3945, signal_3944, signal_3943, signal_1451}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1437 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_3120, signal_3119, signal_3118, signal_1176}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_3948, signal_3947, signal_3946, signal_1452}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1438 ( .a ({signal_3000, signal_2999, signal_2998, signal_1136}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({signal_3951, signal_3950, signal_3949, signal_1453}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1439 ( .a ({signal_2865, signal_2864, signal_2863, signal_1091}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({signal_3954, signal_3953, signal_3952, signal_1454}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1440 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_3063, signal_3062, signal_3061, signal_1157}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({signal_3957, signal_3956, signal_3955, signal_1455}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1441 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_3126, signal_3125, signal_3124, signal_1178}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({signal_3960, signal_3959, signal_3958, signal_1456}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1442 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_3963, signal_3962, signal_3961, signal_1457}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1443 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({signal_3966, signal_3965, signal_3964, signal_1458}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1444 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({signal_3969, signal_3968, signal_3967, signal_1459}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1445 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_3159, signal_3158, signal_3157, signal_1189}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({signal_3972, signal_3971, signal_3970, signal_1460}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1446 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_3162, signal_3161, signal_3160, signal_1190}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({signal_3975, signal_3974, signal_3973, signal_1461}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1447 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_3978, signal_3977, signal_3976, signal_1462}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1448 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_3063, signal_3062, signal_3061, signal_1157}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({signal_3981, signal_3980, signal_3979, signal_1463}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1449 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({signal_3984, signal_3983, signal_3982, signal_1464}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1450 ( .a ({signal_2613, signal_2612, signal_2611, signal_1007}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({signal_3987, signal_3986, signal_3985, signal_1465}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1451 ( .a ({signal_2610, signal_2609, signal_2608, signal_1006}), .b ({signal_3186, signal_3185, signal_3184, signal_1198}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({signal_3990, signal_3989, signal_3988, signal_1466}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1452 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_3027, signal_3026, signal_3025, signal_1145}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_3993, signal_3992, signal_3991, signal_1467}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1453 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_3168, signal_3167, signal_3166, signal_1192}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({signal_3996, signal_3995, signal_3994, signal_1468}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1454 ( .a ({signal_2898, signal_2897, signal_2896, signal_1102}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({signal_3999, signal_3998, signal_3997, signal_1469}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1455 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_3123, signal_3122, signal_3121, signal_1177}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({signal_4002, signal_4001, signal_4000, signal_1470}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1456 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({signal_4005, signal_4004, signal_4003, signal_1471}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1457 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_3165, signal_3164, signal_3163, signal_1191}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_4008, signal_4007, signal_4006, signal_1472}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1458 ( .a ({signal_2640, signal_2639, signal_2638, signal_1016}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({signal_4011, signal_4010, signal_4009, signal_1473}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1459 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_3123, signal_3122, signal_3121, signal_1177}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({signal_4014, signal_4013, signal_4012, signal_1474}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1460 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_3150, signal_3149, signal_3148, signal_1186}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({signal_4017, signal_4016, signal_4015, signal_1475}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1461 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({signal_4020, signal_4019, signal_4018, signal_1476}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1462 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_4023, signal_4022, signal_4021, signal_1477}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1463 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_3210, signal_3209, signal_3208, signal_1206}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({signal_4026, signal_4025, signal_4024, signal_1478}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1464 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({signal_4029, signal_4028, signal_4027, signal_1479}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1465 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_3150, signal_3149, signal_3148, signal_1186}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({signal_4032, signal_4031, signal_4030, signal_1480}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1466 ( .a ({signal_2817, signal_2816, signal_2815, signal_1075}), .b ({signal_2835, signal_2834, signal_2833, signal_1081}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({signal_4035, signal_4034, signal_4033, signal_1481}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1467 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_3096, signal_3095, signal_3094, signal_1168}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_4038, signal_4037, signal_4036, signal_1482}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1468 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_3075, signal_3074, signal_3073, signal_1161}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({signal_4041, signal_4040, signal_4039, signal_1483}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1469 ( .a ({signal_2655, signal_2654, signal_2653, signal_1021}), .b ({signal_2988, signal_2987, signal_2986, signal_1132}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({signal_4044, signal_4043, signal_4042, signal_1484}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1470 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({signal_4047, signal_4046, signal_4045, signal_1485}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1471 ( .a ({signal_2589, signal_2588, signal_2587, signal_999}), .b ({signal_3216, signal_3215, signal_3214, signal_1208}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({signal_4050, signal_4049, signal_4048, signal_1486}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1472 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_4053, signal_4052, signal_4051, signal_1487}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1473 ( .a ({signal_2640, signal_2639, signal_2638, signal_1016}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({signal_4056, signal_4055, signal_4054, signal_1488}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1474 ( .a ({signal_2508, signal_2507, signal_2506, signal_972}), .b ({signal_3195, signal_3194, signal_3193, signal_1201}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({signal_4059, signal_4058, signal_4057, signal_1489}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1475 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_3075, signal_3074, signal_3073, signal_1161}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({signal_4062, signal_4061, signal_4060, signal_1490}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1476 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({signal_4065, signal_4064, signal_4063, signal_1491}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1477 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_3243, signal_3242, signal_3241, signal_1217}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_4068, signal_4067, signal_4066, signal_1492}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1478 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({signal_4071, signal_4070, signal_4069, signal_1493}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1479 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_3159, signal_3158, signal_3157, signal_1189}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({signal_4074, signal_4073, signal_4072, signal_1494}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1480 ( .a ({signal_2520, signal_2519, signal_2518, signal_976}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({signal_4077, signal_4076, signal_4075, signal_1495}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1481 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({signal_4080, signal_4079, signal_4078, signal_1496}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1482 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_4083, signal_4082, signal_4081, signal_1497}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1483 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({signal_4086, signal_4085, signal_4084, signal_1498}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1484 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({signal_4089, signal_4088, signal_4087, signal_1499}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1485 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({signal_4092, signal_4091, signal_4090, signal_1500}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1486 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({signal_4095, signal_4094, signal_4093, signal_1501}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1487 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_4098, signal_4097, signal_4096, signal_1502}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1488 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({signal_4101, signal_4100, signal_4099, signal_1503}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1489 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2949, signal_2948, signal_2947, signal_1119}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({signal_4104, signal_4103, signal_4102, signal_1504}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1490 ( .a ({signal_3690, signal_3689, signal_3688, signal_1366}), .b ({signal_4107, signal_4106, signal_4105, signal_1505}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1491 ( .a ({signal_3693, signal_3692, signal_3691, signal_1367}), .b ({signal_4110, signal_4109, signal_4108, signal_1506}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1497 ( .a ({signal_3711, signal_3710, signal_3709, signal_1373}), .b ({signal_4128, signal_4127, signal_4126, signal_1512}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1498 ( .a ({signal_3714, signal_3713, signal_3712, signal_1374}), .b ({signal_4131, signal_4130, signal_4129, signal_1513}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1502 ( .a ({signal_3726, signal_3725, signal_3724, signal_1378}), .b ({signal_4143, signal_4142, signal_4141, signal_1517}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1503 ( .a ({signal_3729, signal_3728, signal_3727, signal_1379}), .b ({signal_4146, signal_4145, signal_4144, signal_1518}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1508 ( .a ({signal_3747, signal_3746, signal_3745, signal_1385}), .b ({signal_4161, signal_4160, signal_4159, signal_1523}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1509 ( .a ({signal_3750, signal_3749, signal_3748, signal_1386}), .b ({signal_4164, signal_4163, signal_4162, signal_1524}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1510 ( .a ({signal_3753, signal_3752, signal_3751, signal_1387}), .b ({signal_4167, signal_4166, signal_4165, signal_1525}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1511 ( .a ({signal_3756, signal_3755, signal_3754, signal_1388}), .b ({signal_4170, signal_4169, signal_4168, signal_1526}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1512 ( .a ({signal_3759, signal_3758, signal_3757, signal_1389}), .b ({signal_4173, signal_4172, signal_4171, signal_1527}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1514 ( .a ({signal_3768, signal_3767, signal_3766, signal_1392}), .b ({signal_4179, signal_4178, signal_4177, signal_1529}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1515 ( .a ({signal_3771, signal_3770, signal_3769, signal_1393}), .b ({signal_4182, signal_4181, signal_4180, signal_1530}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1516 ( .a ({signal_3774, signal_3773, signal_3772, signal_1394}), .b ({signal_4185, signal_4184, signal_4183, signal_1531}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1517 ( .a ({signal_3777, signal_3776, signal_3775, signal_1395}), .b ({signal_4188, signal_4187, signal_4186, signal_1532}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1518 ( .a ({signal_3780, signal_3779, signal_3778, signal_1396}), .b ({signal_4191, signal_4190, signal_4189, signal_1533}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1519 ( .a ({signal_3783, signal_3782, signal_3781, signal_1397}), .b ({signal_4194, signal_4193, signal_4192, signal_1534}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1521 ( .a ({signal_3789, signal_3788, signal_3787, signal_1399}), .b ({signal_4200, signal_4199, signal_4198, signal_1536}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1522 ( .a ({signal_3792, signal_3791, signal_3790, signal_1400}), .b ({signal_4203, signal_4202, signal_4201, signal_1537}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1523 ( .a ({signal_3795, signal_3794, signal_3793, signal_1401}), .b ({signal_4206, signal_4205, signal_4204, signal_1538}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1524 ( .a ({signal_3798, signal_3797, signal_3796, signal_1402}), .b ({signal_4209, signal_4208, signal_4207, signal_1539}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1525 ( .a ({signal_3801, signal_3800, signal_3799, signal_1403}), .b ({signal_4212, signal_4211, signal_4210, signal_1540}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1526 ( .a ({signal_3804, signal_3803, signal_3802, signal_1404}), .b ({signal_4215, signal_4214, signal_4213, signal_1541}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1527 ( .a ({signal_3807, signal_3806, signal_3805, signal_1405}), .b ({signal_4218, signal_4217, signal_4216, signal_1542}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1528 ( .a ({signal_3810, signal_3809, signal_3808, signal_1406}), .b ({signal_4221, signal_4220, signal_4219, signal_1543}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1529 ( .a ({signal_3813, signal_3812, signal_3811, signal_1407}), .b ({signal_4224, signal_4223, signal_4222, signal_1544}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1530 ( .a ({signal_3816, signal_3815, signal_3814, signal_1408}), .b ({signal_4227, signal_4226, signal_4225, signal_1545}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1531 ( .a ({signal_3819, signal_3818, signal_3817, signal_1409}), .b ({signal_4230, signal_4229, signal_4228, signal_1546}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1534 ( .a ({signal_3828, signal_3827, signal_3826, signal_1412}), .b ({signal_4239, signal_4238, signal_4237, signal_1549}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1535 ( .a ({signal_3831, signal_3830, signal_3829, signal_1413}), .b ({signal_4242, signal_4241, signal_4240, signal_1550}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1536 ( .a ({signal_3834, signal_3833, signal_3832, signal_1414}), .b ({signal_4245, signal_4244, signal_4243, signal_1551}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1537 ( .a ({signal_3837, signal_3836, signal_3835, signal_1415}), .b ({signal_4248, signal_4247, signal_4246, signal_1552}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1540 ( .a ({signal_3849, signal_3848, signal_3847, signal_1419}), .b ({signal_4257, signal_4256, signal_4255, signal_1555}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1541 ( .a ({signal_3852, signal_3851, signal_3850, signal_1420}), .b ({signal_4260, signal_4259, signal_4258, signal_1556}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1542 ( .a ({signal_3855, signal_3854, signal_3853, signal_1421}), .b ({signal_4263, signal_4262, signal_4261, signal_1557}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1545 ( .a ({signal_3864, signal_3863, signal_3862, signal_1424}), .b ({signal_4272, signal_4271, signal_4270, signal_1560}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1546 ( .a ({signal_3867, signal_3866, signal_3865, signal_1425}), .b ({signal_4275, signal_4274, signal_4273, signal_1561}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1547 ( .a ({signal_3870, signal_3869, signal_3868, signal_1426}), .b ({signal_4278, signal_4277, signal_4276, signal_1562}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1548 ( .a ({signal_3873, signal_3872, signal_3871, signal_1427}), .b ({signal_4281, signal_4280, signal_4279, signal_1563}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1549 ( .a ({signal_3876, signal_3875, signal_3874, signal_1428}), .b ({signal_4284, signal_4283, signal_4282, signal_1564}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1550 ( .a ({signal_3879, signal_3878, signal_3877, signal_1429}), .b ({signal_4287, signal_4286, signal_4285, signal_1565}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1551 ( .a ({signal_3882, signal_3881, signal_3880, signal_1430}), .b ({signal_4290, signal_4289, signal_4288, signal_1566}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1552 ( .a ({signal_3885, signal_3884, signal_3883, signal_1431}), .b ({signal_4293, signal_4292, signal_4291, signal_1567}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1553 ( .a ({signal_3888, signal_3887, signal_3886, signal_1432}), .b ({signal_4296, signal_4295, signal_4294, signal_1568}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1554 ( .a ({signal_3891, signal_3890, signal_3889, signal_1433}), .b ({signal_4299, signal_4298, signal_4297, signal_1569}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1555 ( .a ({signal_3894, signal_3893, signal_3892, signal_1434}), .b ({signal_4302, signal_4301, signal_4300, signal_1570}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1556 ( .a ({signal_3897, signal_3896, signal_3895, signal_1435}), .b ({signal_4305, signal_4304, signal_4303, signal_1571}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1557 ( .a ({signal_3900, signal_3899, signal_3898, signal_1436}), .b ({signal_4308, signal_4307, signal_4306, signal_1572}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1558 ( .a ({signal_3903, signal_3902, signal_3901, signal_1437}), .b ({signal_4311, signal_4310, signal_4309, signal_1573}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1559 ( .a ({signal_3906, signal_3905, signal_3904, signal_1438}), .b ({signal_4314, signal_4313, signal_4312, signal_1574}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1560 ( .a ({signal_3909, signal_3908, signal_3907, signal_1439}), .b ({signal_4317, signal_4316, signal_4315, signal_1575}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1561 ( .a ({signal_3912, signal_3911, signal_3910, signal_1440}), .b ({signal_4320, signal_4319, signal_4318, signal_1576}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1562 ( .a ({signal_3915, signal_3914, signal_3913, signal_1441}), .b ({signal_4323, signal_4322, signal_4321, signal_1577}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1563 ( .a ({signal_3918, signal_3917, signal_3916, signal_1442}), .b ({signal_4326, signal_4325, signal_4324, signal_1578}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1564 ( .a ({signal_3921, signal_3920, signal_3919, signal_1443}), .b ({signal_4329, signal_4328, signal_4327, signal_1579}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1565 ( .a ({signal_3924, signal_3923, signal_3922, signal_1444}), .b ({signal_4332, signal_4331, signal_4330, signal_1580}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1566 ( .a ({signal_3927, signal_3926, signal_3925, signal_1445}), .b ({signal_4335, signal_4334, signal_4333, signal_1581}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1567 ( .a ({signal_3933, signal_3932, signal_3931, signal_1447}), .b ({signal_4338, signal_4337, signal_4336, signal_1582}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1568 ( .a ({signal_3936, signal_3935, signal_3934, signal_1448}), .b ({signal_4341, signal_4340, signal_4339, signal_1583}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1569 ( .a ({signal_3939, signal_3938, signal_3937, signal_1449}), .b ({signal_4344, signal_4343, signal_4342, signal_1584}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1570 ( .a ({signal_3942, signal_3941, signal_3940, signal_1450}), .b ({signal_4347, signal_4346, signal_4345, signal_1585}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1571 ( .a ({signal_3945, signal_3944, signal_3943, signal_1451}), .b ({signal_4350, signal_4349, signal_4348, signal_1586}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1572 ( .a ({signal_3948, signal_3947, signal_3946, signal_1452}), .b ({signal_4353, signal_4352, signal_4351, signal_1587}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1573 ( .a ({signal_3951, signal_3950, signal_3949, signal_1453}), .b ({signal_4356, signal_4355, signal_4354, signal_1588}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1574 ( .a ({signal_3954, signal_3953, signal_3952, signal_1454}), .b ({signal_4359, signal_4358, signal_4357, signal_1589}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1575 ( .a ({signal_3957, signal_3956, signal_3955, signal_1455}), .b ({signal_4362, signal_4361, signal_4360, signal_1590}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1576 ( .a ({signal_3960, signal_3959, signal_3958, signal_1456}), .b ({signal_4365, signal_4364, signal_4363, signal_1591}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1577 ( .a ({signal_3963, signal_3962, signal_3961, signal_1457}), .b ({signal_4368, signal_4367, signal_4366, signal_1592}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1578 ( .a ({signal_3966, signal_3965, signal_3964, signal_1458}), .b ({signal_4371, signal_4370, signal_4369, signal_1593}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1579 ( .a ({signal_3969, signal_3968, signal_3967, signal_1459}), .b ({signal_4374, signal_4373, signal_4372, signal_1594}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1580 ( .a ({signal_3972, signal_3971, signal_3970, signal_1460}), .b ({signal_4377, signal_4376, signal_4375, signal_1595}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1581 ( .a ({signal_3978, signal_3977, signal_3976, signal_1462}), .b ({signal_4380, signal_4379, signal_4378, signal_1596}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1582 ( .a ({signal_3981, signal_3980, signal_3979, signal_1463}), .b ({signal_4383, signal_4382, signal_4381, signal_1597}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1583 ( .a ({signal_3984, signal_3983, signal_3982, signal_1464}), .b ({signal_4386, signal_4385, signal_4384, signal_1598}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1584 ( .a ({signal_3987, signal_3986, signal_3985, signal_1465}), .b ({signal_4389, signal_4388, signal_4387, signal_1599}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1585 ( .a ({signal_3990, signal_3989, signal_3988, signal_1466}), .b ({signal_4392, signal_4391, signal_4390, signal_1600}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1586 ( .a ({signal_3993, signal_3992, signal_3991, signal_1467}), .b ({signal_4395, signal_4394, signal_4393, signal_1601}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1587 ( .a ({signal_3996, signal_3995, signal_3994, signal_1468}), .b ({signal_4398, signal_4397, signal_4396, signal_1602}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1588 ( .a ({signal_3999, signal_3998, signal_3997, signal_1469}), .b ({signal_4401, signal_4400, signal_4399, signal_1603}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1589 ( .a ({signal_4002, signal_4001, signal_4000, signal_1470}), .b ({signal_4404, signal_4403, signal_4402, signal_1604}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1590 ( .a ({signal_4005, signal_4004, signal_4003, signal_1471}), .b ({signal_4407, signal_4406, signal_4405, signal_1605}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1591 ( .a ({signal_4008, signal_4007, signal_4006, signal_1472}), .b ({signal_4410, signal_4409, signal_4408, signal_1606}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1592 ( .a ({signal_4011, signal_4010, signal_4009, signal_1473}), .b ({signal_4413, signal_4412, signal_4411, signal_1607}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1593 ( .a ({signal_4014, signal_4013, signal_4012, signal_1474}), .b ({signal_4416, signal_4415, signal_4414, signal_1608}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1594 ( .a ({signal_4017, signal_4016, signal_4015, signal_1475}), .b ({signal_4419, signal_4418, signal_4417, signal_1609}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1595 ( .a ({signal_4020, signal_4019, signal_4018, signal_1476}), .b ({signal_4422, signal_4421, signal_4420, signal_1610}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1596 ( .a ({signal_4023, signal_4022, signal_4021, signal_1477}), .b ({signal_4425, signal_4424, signal_4423, signal_1611}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1597 ( .a ({signal_4029, signal_4028, signal_4027, signal_1479}), .b ({signal_4428, signal_4427, signal_4426, signal_1612}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1598 ( .a ({signal_4032, signal_4031, signal_4030, signal_1480}), .b ({signal_4431, signal_4430, signal_4429, signal_1613}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1599 ( .a ({signal_4035, signal_4034, signal_4033, signal_1481}), .b ({signal_4434, signal_4433, signal_4432, signal_1614}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1600 ( .a ({signal_4038, signal_4037, signal_4036, signal_1482}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1601 ( .a ({signal_4041, signal_4040, signal_4039, signal_1483}), .b ({signal_4440, signal_4439, signal_4438, signal_1616}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1602 ( .a ({signal_4044, signal_4043, signal_4042, signal_1484}), .b ({signal_4443, signal_4442, signal_4441, signal_1617}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1603 ( .a ({signal_4047, signal_4046, signal_4045, signal_1485}), .b ({signal_4446, signal_4445, signal_4444, signal_1618}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1604 ( .a ({signal_4050, signal_4049, signal_4048, signal_1486}), .b ({signal_4449, signal_4448, signal_4447, signal_1619}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1605 ( .a ({signal_4053, signal_4052, signal_4051, signal_1487}), .b ({signal_4452, signal_4451, signal_4450, signal_1620}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1606 ( .a ({signal_4056, signal_4055, signal_4054, signal_1488}), .b ({signal_4455, signal_4454, signal_4453, signal_1621}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1607 ( .a ({signal_4059, signal_4058, signal_4057, signal_1489}), .b ({signal_4458, signal_4457, signal_4456, signal_1622}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1608 ( .a ({signal_4062, signal_4061, signal_4060, signal_1490}), .b ({signal_4461, signal_4460, signal_4459, signal_1623}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1609 ( .a ({signal_4065, signal_4064, signal_4063, signal_1491}), .b ({signal_4464, signal_4463, signal_4462, signal_1624}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1610 ( .a ({signal_4068, signal_4067, signal_4066, signal_1492}), .b ({signal_4467, signal_4466, signal_4465, signal_1625}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1611 ( .a ({signal_4071, signal_4070, signal_4069, signal_1493}), .b ({signal_4470, signal_4469, signal_4468, signal_1626}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1612 ( .a ({signal_4074, signal_4073, signal_4072, signal_1494}), .b ({signal_4473, signal_4472, signal_4471, signal_1627}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1613 ( .a ({signal_4077, signal_4076, signal_4075, signal_1495}), .b ({signal_4476, signal_4475, signal_4474, signal_1628}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1614 ( .a ({signal_4080, signal_4079, signal_4078, signal_1496}), .b ({signal_4479, signal_4478, signal_4477, signal_1629}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1615 ( .a ({signal_4083, signal_4082, signal_4081, signal_1497}), .b ({signal_4482, signal_4481, signal_4480, signal_1630}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1616 ( .a ({signal_4086, signal_4085, signal_4084, signal_1498}), .b ({signal_4485, signal_4484, signal_4483, signal_1631}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1617 ( .a ({signal_4089, signal_4088, signal_4087, signal_1499}), .b ({signal_4488, signal_4487, signal_4486, signal_1632}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1618 ( .a ({signal_4092, signal_4091, signal_4090, signal_1500}), .b ({signal_4491, signal_4490, signal_4489, signal_1633}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1619 ( .a ({signal_4095, signal_4094, signal_4093, signal_1501}), .b ({signal_4494, signal_4493, signal_4492, signal_1634}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1620 ( .a ({signal_4098, signal_4097, signal_4096, signal_1502}), .b ({signal_4497, signal_4496, signal_4495, signal_1635}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1621 ( .a ({signal_4101, signal_4100, signal_4099, signal_1503}), .b ({signal_4500, signal_4499, signal_4498, signal_1636}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1622 ( .a ({signal_4104, signal_4103, signal_4102, signal_1504}), .b ({signal_4503, signal_4502, signal_4501, signal_1637}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1623 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_3282, signal_3281, signal_3280, signal_1230}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({signal_4506, signal_4505, signal_4504, signal_1638}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1624 ( .a ({signal_2763, signal_2762, signal_2761, signal_1057}), .b ({signal_3285, signal_3284, signal_3283, signal_1231}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({signal_4509, signal_4508, signal_4507, signal_1639}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1625 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_3300, signal_3299, signal_3298, signal_1236}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_4512, signal_4511, signal_4510, signal_1640}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1626 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3360, signal_3359, signal_3358, signal_1256}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({signal_4515, signal_4514, signal_4513, signal_1641}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1627 ( .a ({signal_2709, signal_2708, signal_2707, signal_1039}), .b ({signal_3363, signal_3362, signal_3361, signal_1257}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({signal_4518, signal_4517, signal_4516, signal_1642}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1628 ( .a ({signal_2508, signal_2507, signal_2506, signal_972}), .b ({signal_3381, signal_3380, signal_3379, signal_1263}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({signal_4521, signal_4520, signal_4519, signal_1643}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1629 ( .a ({signal_3342, signal_3341, signal_3340, signal_1250}), .b ({signal_3351, signal_3350, signal_3349, signal_1253}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({signal_4524, signal_4523, signal_4522, signal_1644}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1630 ( .a ({signal_3393, signal_3392, signal_3391, signal_1267}), .b ({signal_3396, signal_3395, signal_3394, signal_1268}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_4527, signal_4526, signal_4525, signal_1645}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1631 ( .a ({signal_2730, signal_2729, signal_2728, signal_1046}), .b ({signal_3312, signal_3311, signal_3310, signal_1240}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({signal_4530, signal_4529, signal_4528, signal_1646}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1632 ( .a ({signal_3399, signal_3398, signal_3397, signal_1269}), .b ({signal_3402, signal_3401, signal_3400, signal_1270}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({signal_4533, signal_4532, signal_4531, signal_1647}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1633 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3357, signal_3356, signal_3355, signal_1255}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({signal_4536, signal_4535, signal_4534, signal_1648}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1634 ( .a ({signal_3411, signal_3410, signal_3409, signal_1273}), .b ({signal_3414, signal_3413, signal_3412, signal_1274}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({signal_4539, signal_4538, signal_4537, signal_1649}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1635 ( .a ({signal_2757, signal_2756, signal_2755, signal_1055}), .b ({signal_3354, signal_3353, signal_3352, signal_1254}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_4542, signal_4541, signal_4540, signal_1650}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1636 ( .a ({signal_2520, signal_2519, signal_2518, signal_976}), .b ({signal_3315, signal_3314, signal_3313, signal_1241}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({signal_4545, signal_4544, signal_4543, signal_1651}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1637 ( .a ({signal_3300, signal_3299, signal_3298, signal_1236}), .b ({signal_2769, signal_2768, signal_2767, signal_1059}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({signal_4548, signal_4547, signal_4546, signal_1652}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1638 ( .a ({signal_3432, signal_3431, signal_3430, signal_1280}), .b ({signal_3435, signal_3434, signal_3433, signal_1281}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({signal_4551, signal_4550, signal_4549, signal_1653}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1639 ( .a ({signal_3441, signal_3440, signal_3439, signal_1283}), .b ({signal_3444, signal_3443, signal_3442, signal_1284}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({signal_4554, signal_4553, signal_4552, signal_1654}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1640 ( .a ({signal_3291, signal_3290, signal_3289, signal_1233}), .b ({signal_3450, signal_3449, signal_3448, signal_1286}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_4557, signal_4556, signal_4555, signal_1655}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1641 ( .a ({signal_3303, signal_3302, signal_3301, signal_1237}), .b ({signal_3456, signal_3455, signal_3454, signal_1288}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({signal_4560, signal_4559, signal_4558, signal_1656}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1642 ( .a ({signal_2769, signal_2768, signal_2767, signal_1059}), .b ({signal_3306, signal_3305, signal_3304, signal_1238}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({signal_4563, signal_4562, signal_4561, signal_1657}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1643 ( .a ({signal_3318, signal_3317, signal_3316, signal_1242}), .b ({signal_3321, signal_3320, signal_3319, signal_1243}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({signal_4566, signal_4565, signal_4564, signal_1658}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1645 ( .a ({signal_3474, signal_3473, signal_3472, signal_1294}), .b ({signal_3477, signal_3476, signal_3475, signal_1295}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({signal_4572, signal_4571, signal_4570, signal_1660}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1646 ( .a ({signal_3306, signal_3305, signal_3304, signal_1238}), .b ({signal_3498, signal_3497, signal_3496, signal_1302}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_4575, signal_4574, signal_4573, signal_1661}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1647 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_3510, signal_3509, signal_3508, signal_1306}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({signal_4578, signal_4577, signal_4576, signal_1662}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1648 ( .a ({signal_3348, signal_3347, signal_3346, signal_1252}), .b ({signal_3522, signal_3521, signal_3520, signal_1310}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({signal_4581, signal_4580, signal_4579, signal_1663}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1649 ( .a ({signal_2715, signal_2714, signal_2713, signal_1041}), .b ({signal_3741, signal_3740, signal_3739, signal_1383}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({signal_4584, signal_4583, signal_4582, signal_1664}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1650 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({signal_4587, signal_4586, signal_4585, signal_1665}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1651 ( .a ({signal_3324, signal_3323, signal_3322, signal_1244}), .b ({signal_3525, signal_3524, signal_3523, signal_1311}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_4590, signal_4589, signal_4588, signal_1666}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1653 ( .a ({signal_3720, signal_3719, signal_3718, signal_1376}), .b ({signal_3543, signal_3542, signal_3541, signal_1317}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({signal_4596, signal_4595, signal_4594, signal_1668}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1654 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3549, signal_3548, signal_3547, signal_1319}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({signal_4599, signal_4598, signal_4597, signal_1669}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1655 ( .a ({signal_3762, signal_3761, signal_3760, signal_1390}), .b ({signal_2787, signal_2786, signal_2785, signal_1065}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({signal_4602, signal_4601, signal_4600, signal_1670}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1656 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({signal_4605, signal_4604, signal_4603, signal_1671}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1657 ( .a ({signal_3372, signal_3371, signal_3370, signal_1260}), .b ({signal_3492, signal_3491, signal_3490, signal_1300}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_4608, signal_4607, signal_4606, signal_1672}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1658 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_3555, signal_3554, signal_3553, signal_1321}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({signal_4611, signal_4610, signal_4609, signal_1673}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1659 ( .a ({signal_3540, signal_3539, signal_3538, signal_1316}), .b ({signal_3558, signal_3557, signal_3556, signal_1322}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({signal_4614, signal_4613, signal_4612, signal_1674}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1660 ( .a ({signal_2781, signal_2780, signal_2779, signal_1063}), .b ({signal_3561, signal_3560, signal_3559, signal_1323}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({signal_4617, signal_4616, signal_4615, signal_1675}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1661 ( .a ({signal_3564, signal_3563, signal_3562, signal_1324}), .b ({signal_3567, signal_3566, signal_3565, signal_1325}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({signal_4620, signal_4619, signal_4618, signal_1676}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1663 ( .a ({signal_3312, signal_3311, signal_3310, signal_1240}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_4626, signal_4625, signal_4624, signal_1678}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1664 ( .a ({signal_3384, signal_3383, signal_3382, signal_1264}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({signal_4629, signal_4628, signal_4627, signal_1679}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1665 ( .a ({signal_3318, signal_3317, signal_3316, signal_1242}), .b ({signal_3588, signal_3587, signal_3586, signal_1332}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({signal_4632, signal_4631, signal_4630, signal_1680}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1666 ( .a ({signal_3390, signal_3389, signal_3388, signal_1266}), .b ({signal_3594, signal_3593, signal_3592, signal_1334}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({signal_4635, signal_4634, signal_4633, signal_1681}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1667 ( .a ({signal_3483, signal_3482, signal_3481, signal_1297}), .b ({signal_3603, signal_3602, signal_3601, signal_1337}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({signal_4638, signal_4637, signal_4636, signal_1682}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1668 ( .a ({signal_3405, signal_3404, signal_3403, signal_1271}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_4641, signal_4640, signal_4639, signal_1683}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1669 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({signal_4644, signal_4643, signal_4642, signal_1684}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1670 ( .a ({signal_3459, signal_3458, signal_3457, signal_1289}), .b ({signal_3612, signal_3611, signal_3610, signal_1340}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({signal_4647, signal_4646, signal_4645, signal_1685}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1671 ( .a ({signal_2694, signal_2693, signal_2692, signal_1034}), .b ({signal_3615, signal_3614, signal_3613, signal_1341}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({signal_4650, signal_4649, signal_4648, signal_1686}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1673 ( .a ({signal_3420, signal_3419, signal_3418, signal_1276}), .b ({signal_3582, signal_3581, signal_3580, signal_1330}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({signal_4656, signal_4655, signal_4654, signal_1688}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1674 ( .a ({signal_3546, signal_3545, signal_3544, signal_1318}), .b ({signal_3846, signal_3845, signal_3844, signal_1418}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_4659, signal_4658, signal_4657, signal_1689}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1675 ( .a ({signal_3369, signal_3368, signal_3367, signal_1259}), .b ({signal_3564, signal_3563, signal_3562, signal_1324}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({signal_4662, signal_4661, signal_4660, signal_1690}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1676 ( .a ({signal_3423, signal_3422, signal_3421, signal_1277}), .b ({signal_3630, signal_3629, signal_3628, signal_1346}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({signal_4665, signal_4664, signal_4663, signal_1691}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1677 ( .a ({signal_3633, signal_3632, signal_3631, signal_1347}), .b ({signal_3636, signal_3635, signal_3634, signal_1348}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({signal_4668, signal_4667, signal_4666, signal_1692}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1678 ( .a ({signal_3342, signal_3341, signal_3340, signal_1250}), .b ({signal_3639, signal_3638, signal_3637, signal_1349}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({signal_4671, signal_4670, signal_4669, signal_1693}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1679 ( .a ({signal_3645, signal_3644, signal_3643, signal_1351}), .b ({signal_3648, signal_3647, signal_3646, signal_1352}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_4674, signal_4673, signal_4672, signal_1694}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1680 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3519, signal_3518, signal_3517, signal_1309}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({signal_4677, signal_4676, signal_4675, signal_1695}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1681 ( .a ({signal_3657, signal_3656, signal_3655, signal_1355}), .b ({signal_3660, signal_3659, signal_3658, signal_1356}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({signal_4680, signal_4679, signal_4678, signal_1696}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1682 ( .a ({signal_3537, signal_3536, signal_3535, signal_1315}), .b ({signal_3663, signal_3662, signal_3661, signal_1357}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({signal_4683, signal_4682, signal_4681, signal_1697}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1684 ( .a ({signal_3459, signal_3458, signal_3457, signal_1289}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({signal_4689, signal_4688, signal_4687, signal_1699}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1687 ( .a ({signal_3321, signal_3320, signal_3319, signal_1243}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_4698, signal_4697, signal_4696, signal_1702}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1693 ( .a ({signal_3462, signal_3461, signal_3460, signal_1290}), .b ({signal_3507, signal_3506, signal_3505, signal_1305}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({signal_4716, signal_4715, signal_4714, signal_1708}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1698 ( .a ({signal_3471, signal_3470, signal_3469, signal_1293}), .b ({signal_3684, signal_3683, signal_3682, signal_1364}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({signal_4731, signal_4730, signal_4729, signal_1713}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1700 ( .a ({signal_4506, signal_4505, signal_4504, signal_1638}), .b ({signal_4737, signal_4736, signal_4735, signal_1715}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1701 ( .a ({signal_4509, signal_4508, signal_4507, signal_1639}), .b ({signal_4740, signal_4739, signal_4738, signal_1716}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1702 ( .a ({signal_4515, signal_4514, signal_4513, signal_1641}), .b ({signal_4743, signal_4742, signal_4741, signal_1717}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1703 ( .a ({signal_4518, signal_4517, signal_4516, signal_1642}), .b ({signal_4746, signal_4745, signal_4744, signal_1718}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1704 ( .a ({signal_4521, signal_4520, signal_4519, signal_1643}), .b ({signal_4749, signal_4748, signal_4747, signal_1719}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1705 ( .a ({signal_4524, signal_4523, signal_4522, signal_1644}), .b ({signal_4752, signal_4751, signal_4750, signal_1720}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1706 ( .a ({signal_4530, signal_4529, signal_4528, signal_1646}), .b ({signal_4755, signal_4754, signal_4753, signal_1721}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1707 ( .a ({signal_4533, signal_4532, signal_4531, signal_1647}), .b ({signal_4758, signal_4757, signal_4756, signal_1722}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1708 ( .a ({signal_4536, signal_4535, signal_4534, signal_1648}), .b ({signal_4761, signal_4760, signal_4759, signal_1723}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1709 ( .a ({signal_4542, signal_4541, signal_4540, signal_1650}), .b ({signal_4764, signal_4763, signal_4762, signal_1724}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1710 ( .a ({signal_4545, signal_4544, signal_4543, signal_1651}), .b ({signal_4767, signal_4766, signal_4765, signal_1725}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1711 ( .a ({signal_4548, signal_4547, signal_4546, signal_1652}), .b ({signal_4770, signal_4769, signal_4768, signal_1726}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1712 ( .a ({signal_4560, signal_4559, signal_4558, signal_1656}), .b ({signal_4773, signal_4772, signal_4771, signal_1727}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1713 ( .a ({signal_4563, signal_4562, signal_4561, signal_1657}), .b ({signal_4776, signal_4775, signal_4774, signal_1728}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1714 ( .a ({signal_4566, signal_4565, signal_4564, signal_1658}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1716 ( .a ({signal_4578, signal_4577, signal_4576, signal_1662}), .b ({signal_4785, signal_4784, signal_4783, signal_1731}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1717 ( .a ({signal_4581, signal_4580, signal_4579, signal_1663}), .b ({signal_4788, signal_4787, signal_4786, signal_1732}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1718 ( .a ({signal_4584, signal_4583, signal_4582, signal_1664}), .b ({signal_4791, signal_4790, signal_4789, signal_1733}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1719 ( .a ({signal_4587, signal_4586, signal_4585, signal_1665}), .b ({signal_4794, signal_4793, signal_4792, signal_1734}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1720 ( .a ({signal_4590, signal_4589, signal_4588, signal_1666}), .b ({signal_4797, signal_4796, signal_4795, signal_1735}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1722 ( .a ({signal_4599, signal_4598, signal_4597, signal_1669}), .b ({signal_4803, signal_4802, signal_4801, signal_1737}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1723 ( .a ({signal_4611, signal_4610, signal_4609, signal_1673}), .b ({signal_4806, signal_4805, signal_4804, signal_1738}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1724 ( .a ({signal_4620, signal_4619, signal_4618, signal_1676}), .b ({signal_4809, signal_4808, signal_4807, signal_1739}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1726 ( .a ({signal_4626, signal_4625, signal_4624, signal_1678}), .b ({signal_4815, signal_4814, signal_4813, signal_1741}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1727 ( .a ({signal_4629, signal_4628, signal_4627, signal_1679}), .b ({signal_4818, signal_4817, signal_4816, signal_1742}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1728 ( .a ({signal_4632, signal_4631, signal_4630, signal_1680}), .b ({signal_4821, signal_4820, signal_4819, signal_1743}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1729 ( .a ({signal_4635, signal_4634, signal_4633, signal_1681}), .b ({signal_4824, signal_4823, signal_4822, signal_1744}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1730 ( .a ({signal_4638, signal_4637, signal_4636, signal_1682}), .b ({signal_4827, signal_4826, signal_4825, signal_1745}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1731 ( .a ({signal_4650, signal_4649, signal_4648, signal_1686}), .b ({signal_4830, signal_4829, signal_4828, signal_1746}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1732 ( .a ({signal_4659, signal_4658, signal_4657, signal_1689}), .b ({signal_4833, signal_4832, signal_4831, signal_1747}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1733 ( .a ({signal_4671, signal_4670, signal_4669, signal_1693}), .b ({signal_4836, signal_4835, signal_4834, signal_1748}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1734 ( .a ({signal_4680, signal_4679, signal_4678, signal_1696}), .b ({signal_4839, signal_4838, signal_4837, signal_1749}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1735 ( .a ({signal_4683, signal_4682, signal_4681, signal_1697}), .b ({signal_4842, signal_4841, signal_4840, signal_1750}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1736 ( .a ({signal_4689, signal_4688, signal_4687, signal_1699}), .b ({signal_4845, signal_4844, signal_4843, signal_1751}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1739 ( .a ({signal_4698, signal_4697, signal_4696, signal_1702}), .b ({signal_4854, signal_4853, signal_4852, signal_1754}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1745 ( .a ({signal_4716, signal_4715, signal_4714, signal_1708}), .b ({signal_4872, signal_4871, signal_4870, signal_1760}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1749 ( .a ({signal_4731, signal_4730, signal_4729, signal_1713}), .b ({signal_4884, signal_4883, signal_4882, signal_1764}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1751 ( .a ({signal_2898, signal_2897, signal_2896, signal_1102}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({signal_4890, signal_4889, signal_4888, signal_1766}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1753 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({signal_4116, signal_4115, signal_4114, signal_1508}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({signal_4896, signal_4895, signal_4894, signal_1768}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1754 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_4119, signal_4118, signal_4117, signal_1509}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_4899, signal_4898, signal_4897, signal_1769}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1755 ( .a ({signal_2841, signal_2840, signal_2839, signal_1083}), .b ({signal_4122, signal_4121, signal_4120, signal_1510}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({signal_4902, signal_4901, signal_4900, signal_1770}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1756 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({signal_4905, signal_4904, signal_4903, signal_1771}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1757 ( .a ({signal_2988, signal_2987, signal_2986, signal_1132}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({signal_4908, signal_4907, signal_4906, signal_1772}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1758 ( .a ({signal_2589, signal_2588, signal_2587, signal_999}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({signal_4911, signal_4910, signal_4909, signal_1773}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1760 ( .a ({signal_2580, signal_2579, signal_2578, signal_996}), .b ({signal_4134, signal_4133, signal_4132, signal_1514}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_4917, signal_4916, signal_4915, signal_1775}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1761 ( .a ({signal_2574, signal_2573, signal_2572, signal_994}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}), .clk ( clk ), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({signal_4920, signal_4919, signal_4918, signal_1776}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1762 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_4140, signal_4139, signal_4138, signal_1516}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({signal_4923, signal_4922, signal_4921, signal_1777}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1764 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_4149, signal_4148, signal_4147, signal_1519}), .clk ( clk ), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({signal_4929, signal_4928, signal_4927, signal_1779}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1765 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({signal_4932, signal_4931, signal_4930, signal_1780}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1766 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}), .clk ( clk ), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_4935, signal_4934, signal_4933, signal_1781}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1767 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}), .clk ( clk ), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({signal_4938, signal_4937, signal_4936, signal_1782}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1769 ( .a ({signal_2826, signal_2825, signal_2824, signal_1078}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}), .clk ( clk ), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({signal_4944, signal_4943, signal_4942, signal_1784}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1770 ( .a ({signal_2847, signal_2846, signal_2845, signal_1085}), .b ({signal_4176, signal_4175, signal_4174, signal_1528}), .clk ( clk ), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({signal_4947, signal_4946, signal_4945, signal_1785}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1772 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({signal_4953, signal_4952, signal_4951, signal_1787}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1773 ( .a ({signal_3051, signal_3050, signal_3049, signal_1153}), .b ({signal_4197, signal_4196, signal_4195, signal_1535}), .clk ( clk ), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_4956, signal_4955, signal_4954, signal_1788}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1776 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}), .clk ( clk ), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({signal_4965, signal_4964, signal_4963, signal_1791}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1778 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_4233, signal_4232, signal_4231, signal_1547}), .clk ( clk ), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({signal_4971, signal_4970, signal_4969, signal_1793}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1779 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_4236, signal_4235, signal_4234, signal_1548}), .clk ( clk ), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({signal_4974, signal_4973, signal_4972, signal_1794}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1782 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_4251, signal_4250, signal_4249, signal_1553}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({signal_4983, signal_4982, signal_4981, signal_1797}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1783 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_4254, signal_4253, signal_4252, signal_1554}), .clk ( clk ), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_4986, signal_4985, signal_4984, signal_1798}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1784 ( .a ({signal_2838, signal_2837, signal_2836, signal_1082}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}), .clk ( clk ), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({signal_4989, signal_4988, signal_4987, signal_1799}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1785 ( .a ({signal_2613, signal_2612, signal_2611, signal_1007}), .b ({signal_4266, signal_4265, signal_4264, signal_1558}), .clk ( clk ), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({signal_4992, signal_4991, signal_4990, signal_1800}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1786 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_4269, signal_4268, signal_4267, signal_1559}), .clk ( clk ), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({signal_4995, signal_4994, signal_4993, signal_1801}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1835 ( .a ({signal_4890, signal_4889, signal_4888, signal_1766}), .b ({signal_5142, signal_5141, signal_5140, signal_1850}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1836 ( .a ({signal_4902, signal_4901, signal_4900, signal_1770}), .b ({signal_5145, signal_5144, signal_5143, signal_1851}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1837 ( .a ({signal_4908, signal_4907, signal_4906, signal_1772}), .b ({signal_5148, signal_5147, signal_5146, signal_1852}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1838 ( .a ({signal_4911, signal_4910, signal_4909, signal_1773}), .b ({signal_5151, signal_5150, signal_5149, signal_1853}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1839 ( .a ({signal_4917, signal_4916, signal_4915, signal_1775}), .b ({signal_5154, signal_5153, signal_5152, signal_1854}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1840 ( .a ({signal_4920, signal_4919, signal_4918, signal_1776}), .b ({signal_5157, signal_5156, signal_5155, signal_1855}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1841 ( .a ({signal_4923, signal_4922, signal_4921, signal_1777}), .b ({signal_5160, signal_5159, signal_5158, signal_1856}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1843 ( .a ({signal_4929, signal_4928, signal_4927, signal_1779}), .b ({signal_5166, signal_5165, signal_5164, signal_1858}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1844 ( .a ({signal_4932, signal_4931, signal_4930, signal_1780}), .b ({signal_5169, signal_5168, signal_5167, signal_1859}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1845 ( .a ({signal_4935, signal_4934, signal_4933, signal_1781}), .b ({signal_5172, signal_5171, signal_5170, signal_1860}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1846 ( .a ({signal_4944, signal_4943, signal_4942, signal_1784}), .b ({signal_5175, signal_5174, signal_5173, signal_1861}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1847 ( .a ({signal_4947, signal_4946, signal_4945, signal_1785}), .b ({signal_5178, signal_5177, signal_5176, signal_1862}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1848 ( .a ({signal_4953, signal_4952, signal_4951, signal_1787}), .b ({signal_5181, signal_5180, signal_5179, signal_1863}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1849 ( .a ({signal_4956, signal_4955, signal_4954, signal_1788}), .b ({signal_5184, signal_5183, signal_5182, signal_1864}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1850 ( .a ({signal_4965, signal_4964, signal_4963, signal_1791}), .b ({signal_5187, signal_5186, signal_5185, signal_1865}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1851 ( .a ({signal_4971, signal_4970, signal_4969, signal_1793}), .b ({signal_5190, signal_5189, signal_5188, signal_1866}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1852 ( .a ({signal_4974, signal_4973, signal_4972, signal_1794}), .b ({signal_5193, signal_5192, signal_5191, signal_1867}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1854 ( .a ({signal_4983, signal_4982, signal_4981, signal_1797}), .b ({signal_5199, signal_5198, signal_5197, signal_1869}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1855 ( .a ({signal_4986, signal_4985, signal_4984, signal_1798}), .b ({signal_5202, signal_5201, signal_5200, signal_1870}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1856 ( .a ({signal_4989, signal_4988, signal_4987, signal_1799}), .b ({signal_5205, signal_5204, signal_5203, signal_1871}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1857 ( .a ({signal_4992, signal_4991, signal_4990, signal_1800}), .b ({signal_5208, signal_5207, signal_5206, signal_1872}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1858 ( .a ({signal_4995, signal_4994, signal_4993, signal_1801}), .b ({signal_5211, signal_5210, signal_5209, signal_1873}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1644 ( .a ({signal_3468, signal_3467, signal_3466, signal_1292}), .b ({signal_3471, signal_3470, signal_3469, signal_1293}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({signal_4569, signal_4568, signal_4567, signal_1659}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1652 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_3747, signal_3746, signal_3745, signal_1385}), .clk ( clk ), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_4593, signal_4592, signal_4591, signal_1667}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1662 ( .a ({signal_3576, signal_3575, signal_3574, signal_1328}), .b ({signal_3579, signal_3578, signal_3577, signal_1329}), .clk ( clk ), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({signal_4623, signal_4622, signal_4621, signal_1677}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1672 ( .a ({signal_3618, signal_3617, signal_3616, signal_1342}), .b ({signal_3621, signal_3620, signal_3619, signal_1343}), .clk ( clk ), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({signal_4653, signal_4652, signal_4651, signal_1687}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1683 ( .a ({signal_3438, signal_3437, signal_3436, signal_1282}), .b ({signal_3666, signal_3665, signal_3664, signal_1358}), .clk ( clk ), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({signal_4686, signal_4685, signal_4684, signal_1698}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1685 ( .a ({signal_3465, signal_3464, signal_3463, signal_1291}), .b ({signal_3672, signal_3671, signal_3670, signal_1360}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({signal_4692, signal_4691, signal_4690, signal_1700}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1686 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_3930, signal_3929, signal_3928, signal_1446}), .clk ( clk ), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_4695, signal_4694, signal_4693, signal_1701}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1688 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_3930, signal_3929, signal_3928, signal_1446}), .clk ( clk ), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({signal_4701, signal_4700, signal_4699, signal_1703}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1689 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_3972, signal_3971, signal_3970, signal_1460}), .clk ( clk ), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({signal_4704, signal_4703, signal_4702, signal_1704}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1690 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_3975, signal_3974, signal_3973, signal_1461}), .clk ( clk ), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({signal_4707, signal_4706, signal_4705, signal_1705}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1691 ( .a ({signal_2520, signal_2519, signal_2518, signal_976}), .b ({signal_3978, signal_3977, signal_3976, signal_1462}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({signal_4710, signal_4709, signal_4708, signal_1706}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1692 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_3942, signal_3941, signal_3940, signal_1450}), .clk ( clk ), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_4713, signal_4712, signal_4711, signal_1707}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1694 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_4026, signal_4025, signal_4024, signal_1478}), .clk ( clk ), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({signal_4719, signal_4718, signal_4717, signal_1709}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1695 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_3681, signal_3680, signal_3679, signal_1363}), .clk ( clk ), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({signal_4722, signal_4721, signal_4720, signal_1710}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1696 ( .a ({signal_2730, signal_2729, signal_2728, signal_1046}), .b ({signal_3897, signal_3896, signal_3895, signal_1435}), .clk ( clk ), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({signal_4725, signal_4724, signal_4723, signal_1711}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1697 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_4014, signal_4013, signal_4012, signal_1474}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({signal_4728, signal_4727, signal_4726, signal_1712}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1699 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_4083, signal_4082, signal_4081, signal_1497}), .clk ( clk ), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_4734, signal_4733, signal_4732, signal_1714}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1715 ( .a ({signal_4569, signal_4568, signal_4567, signal_1659}), .b ({signal_4782, signal_4781, signal_4780, signal_1730}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1721 ( .a ({signal_4593, signal_4592, signal_4591, signal_1667}), .b ({signal_4800, signal_4799, signal_4798, signal_1736}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1725 ( .a ({signal_4623, signal_4622, signal_4621, signal_1677}), .b ({signal_4812, signal_4811, signal_4810, signal_1740}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1737 ( .a ({signal_4692, signal_4691, signal_4690, signal_1700}), .b ({signal_4848, signal_4847, signal_4846, signal_1752}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1738 ( .a ({signal_4695, signal_4694, signal_4693, signal_1701}), .b ({signal_4851, signal_4850, signal_4849, signal_1753}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1740 ( .a ({signal_4701, signal_4700, signal_4699, signal_1703}), .b ({signal_4857, signal_4856, signal_4855, signal_1755}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1741 ( .a ({signal_4704, signal_4703, signal_4702, signal_1704}), .b ({signal_4860, signal_4859, signal_4858, signal_1756}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1742 ( .a ({signal_4707, signal_4706, signal_4705, signal_1705}), .b ({signal_4863, signal_4862, signal_4861, signal_1757}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1743 ( .a ({signal_4710, signal_4709, signal_4708, signal_1706}), .b ({signal_4866, signal_4865, signal_4864, signal_1758}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1744 ( .a ({signal_4713, signal_4712, signal_4711, signal_1707}), .b ({signal_4869, signal_4868, signal_4867, signal_1759}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1746 ( .a ({signal_4719, signal_4718, signal_4717, signal_1709}), .b ({signal_4875, signal_4874, signal_4873, signal_1761}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1747 ( .a ({signal_4725, signal_4724, signal_4723, signal_1711}), .b ({signal_4878, signal_4877, signal_4876, signal_1762}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1748 ( .a ({signal_4728, signal_4727, signal_4726, signal_1712}), .b ({signal_4881, signal_4880, signal_4879, signal_1763}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1750 ( .a ({signal_4734, signal_4733, signal_4732, signal_1714}), .b ({signal_4887, signal_4886, signal_4885, signal_1765}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1752 ( .a ({signal_4185, signal_4184, signal_4183, signal_1531}), .b ({signal_4188, signal_4187, signal_4186, signal_1532}), .clk ( clk ), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({signal_4893, signal_4892, signal_4891, signal_1767}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1759 ( .a ({signal_2736, signal_2735, signal_2734, signal_1048}), .b ({signal_4128, signal_4127, signal_4126, signal_1512}), .clk ( clk ), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({signal_4914, signal_4913, signal_4912, signal_1774}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1763 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_4143, signal_4142, signal_4141, signal_1517}), .clk ( clk ), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({signal_4926, signal_4925, signal_4924, signal_1778}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1768 ( .a ({signal_4167, signal_4166, signal_4165, signal_1525}), .b ({signal_4170, signal_4169, signal_4168, signal_1526}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({signal_4941, signal_4940, signal_4939, signal_1783}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1771 ( .a ({signal_4161, signal_4160, signal_4159, signal_1523}), .b ({signal_4182, signal_4181, signal_4180, signal_1530}), .clk ( clk ), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_4950, signal_4949, signal_4948, signal_1786}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1774 ( .a ({signal_3378, signal_3377, signal_3376, signal_1262}), .b ({signal_4200, signal_4199, signal_4198, signal_1536}), .clk ( clk ), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({signal_4959, signal_4958, signal_4957, signal_1789}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1775 ( .a ({signal_4215, signal_4214, signal_4213, signal_1541}), .b ({signal_4218, signal_4217, signal_4216, signal_1542}), .clk ( clk ), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({signal_4962, signal_4961, signal_4960, signal_1790}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1777 ( .a ({signal_3324, signal_3323, signal_3322, signal_1244}), .b ({signal_4230, signal_4229, signal_4228, signal_1546}), .clk ( clk ), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({signal_4968, signal_4967, signal_4966, signal_1792}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1780 ( .a ({signal_3417, signal_3416, signal_3415, signal_1275}), .b ({signal_4539, signal_4538, signal_4537, signal_1649}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({signal_4977, signal_4976, signal_4975, signal_1795}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1781 ( .a ({signal_4374, signal_4373, signal_4372, signal_1594}), .b ({signal_4425, signal_4424, signal_4423, signal_1611}), .clk ( clk ), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_4980, signal_4979, signal_4978, signal_1796}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1787 ( .a ({signal_3357, signal_3356, signal_3355, signal_1255}), .b ({signal_4275, signal_4274, signal_4273, signal_1561}), .clk ( clk ), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({signal_4998, signal_4997, signal_4996, signal_1802}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1788 ( .a ({signal_4281, signal_4280, signal_4279, signal_1563}), .b ({signal_3651, signal_3650, signal_3649, signal_1353}), .clk ( clk ), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({signal_5001, signal_5000, signal_4999, signal_1803}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1789 ( .a ({signal_3639, signal_3638, signal_3637, signal_1349}), .b ({signal_4551, signal_4550, signal_4549, signal_1653}), .clk ( clk ), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({signal_5004, signal_5003, signal_5002, signal_1804}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1790 ( .a ({signal_3288, signal_3287, signal_3286, signal_1232}), .b ({signal_4554, signal_4553, signal_4552, signal_1654}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({signal_5007, signal_5006, signal_5005, signal_1805}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1791 ( .a ({signal_3447, signal_3446, signal_3445, signal_1285}), .b ({signal_4557, signal_4556, signal_4555, signal_1655}), .clk ( clk ), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_5010, signal_5009, signal_5008, signal_1806}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1792 ( .a ({signal_4290, signal_4289, signal_4288, signal_1566}), .b ({signal_4293, signal_4292, signal_4291, signal_1567}), .clk ( clk ), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({signal_5013, signal_5012, signal_5011, signal_1807}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1793 ( .a ({signal_3453, signal_3452, signal_3451, signal_1287}), .b ({signal_4296, signal_4295, signal_4294, signal_1568}), .clk ( clk ), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({signal_5016, signal_5015, signal_5014, signal_1808}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1794 ( .a ({signal_4512, signal_4511, signal_4510, signal_1640}), .b ({signal_4299, signal_4298, signal_4297, signal_1569}), .clk ( clk ), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({signal_5019, signal_5018, signal_5017, signal_1809}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1795 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_4305, signal_4304, signal_4303, signal_1571}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({signal_5022, signal_5021, signal_5020, signal_1810}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1796 ( .a ({signal_4131, signal_4130, signal_4129, signal_1513}), .b ({signal_4308, signal_4307, signal_4306, signal_1572}), .clk ( clk ), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_5025, signal_5024, signal_5023, signal_1811}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1797 ( .a ({signal_3327, signal_3326, signal_3325, signal_1245}), .b ({signal_4311, signal_4310, signal_4309, signal_1573}), .clk ( clk ), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({signal_5028, signal_5027, signal_5026, signal_1812}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1798 ( .a ({signal_3330, signal_3329, signal_3328, signal_1246}), .b ({signal_4572, signal_4571, signal_4570, signal_1660}), .clk ( clk ), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({signal_5031, signal_5030, signal_5029, signal_1813}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1799 ( .a ({signal_2781, signal_2780, signal_2779, signal_1063}), .b ({signal_4314, signal_4313, signal_4312, signal_1574}), .clk ( clk ), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({signal_5034, signal_5033, signal_5032, signal_1814}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1800 ( .a ({signal_3495, signal_3494, signal_3493, signal_1301}), .b ({signal_4323, signal_4322, signal_4321, signal_1577}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({signal_5037, signal_5036, signal_5035, signal_1815}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1801 ( .a ({signal_3339, signal_3338, signal_3337, signal_1249}), .b ({signal_4575, signal_4574, signal_4573, signal_1661}), .clk ( clk ), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_5040, signal_5039, signal_5038, signal_1816}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1802 ( .a ({signal_3501, signal_3500, signal_3499, signal_1303}), .b ({signal_4290, signal_4289, signal_4288, signal_1566}), .clk ( clk ), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({signal_5043, signal_5042, signal_5041, signal_1817}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1803 ( .a ({signal_4329, signal_4328, signal_4327, signal_1579}), .b ({signal_4332, signal_4331, signal_4330, signal_1580}), .clk ( clk ), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({signal_5046, signal_5045, signal_5044, signal_1818}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1804 ( .a ({signal_4164, signal_4163, signal_4162, signal_1524}), .b ({signal_4347, signal_4346, signal_4345, signal_1585}), .clk ( clk ), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({signal_5049, signal_5048, signal_5047, signal_1819}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1805 ( .a ({signal_4314, signal_4313, signal_4312, signal_1574}), .b ({signal_4350, signal_4349, signal_4348, signal_1586}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({signal_5052, signal_5051, signal_5050, signal_1820}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1806 ( .a ({signal_2754, signal_2753, signal_2752, signal_1054}), .b ({signal_4596, signal_4595, signal_4594, signal_1668}), .clk ( clk ), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_5055, signal_5054, signal_5053, signal_1821}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1807 ( .a ({signal_3351, signal_3350, signal_3349, signal_1253}), .b ({signal_4590, signal_4589, signal_4588, signal_1666}), .clk ( clk ), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({signal_5058, signal_5057, signal_5056, signal_1822}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1808 ( .a ({signal_3369, signal_3368, signal_3367, signal_1259}), .b ({signal_4602, signal_4601, signal_4600, signal_1670}), .clk ( clk ), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({signal_5061, signal_5060, signal_5059, signal_1823}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1809 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_4605, signal_4604, signal_4603, signal_1671}), .clk ( clk ), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({signal_5064, signal_5063, signal_5062, signal_1824}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1810 ( .a ({signal_4479, signal_4478, signal_4477, signal_1629}), .b ({signal_4482, signal_4481, signal_4480, signal_1630}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({signal_5067, signal_5066, signal_5065, signal_1825}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1811 ( .a ({signal_4179, signal_4178, signal_4177, signal_1529}), .b ({signal_4608, signal_4607, signal_4606, signal_1672}), .clk ( clk ), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_5070, signal_5069, signal_5068, signal_1826}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1812 ( .a ({signal_4206, signal_4205, signal_4204, signal_1538}), .b ({signal_4389, signal_4388, signal_4387, signal_1599}), .clk ( clk ), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({signal_5073, signal_5072, signal_5071, signal_1827}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1813 ( .a ({signal_4224, signal_4223, signal_4222, signal_1544}), .b ({signal_4407, signal_4406, signal_4405, signal_1605}), .clk ( clk ), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({signal_5076, signal_5075, signal_5074, signal_1828}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1814 ( .a ({signal_4227, signal_4226, signal_4225, signal_1545}), .b ({signal_4413, signal_4412, signal_4411, signal_1607}), .clk ( clk ), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({signal_5079, signal_5078, signal_5077, signal_1829}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1815 ( .a ({signal_3609, signal_3608, signal_3607, signal_1339}), .b ({signal_4416, signal_4415, signal_4414, signal_1608}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({signal_5082, signal_5081, signal_5080, signal_1830}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1816 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_4644, signal_4643, signal_4642, signal_1684}), .clk ( clk ), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_5085, signal_5084, signal_5083, signal_1831}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1817 ( .a ({signal_3408, signal_3407, signal_3406, signal_1272}), .b ({signal_4647, signal_4646, signal_4645, signal_1685}), .clk ( clk ), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({signal_5088, signal_5087, signal_5086, signal_1832}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1818 ( .a ({signal_4305, signal_4304, signal_4303, signal_1571}), .b ({signal_4380, signal_4379, signal_4378, signal_1596}), .clk ( clk ), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({signal_5091, signal_5090, signal_5089, signal_1833}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1820 ( .a ({signal_3624, signal_3623, signal_3622, signal_1344}), .b ({signal_4422, signal_4421, signal_4420, signal_1610}), .clk ( clk ), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({signal_5097, signal_5096, signal_5095, signal_1835}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1821 ( .a ({signal_2778, signal_2777, signal_2776, signal_1062}), .b ({signal_4428, signal_4427, signal_4426, signal_1612}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({signal_5100, signal_5099, signal_5098, signal_1836}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1822 ( .a ({signal_3627, signal_3626, signal_3625, signal_1345}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}), .clk ( clk ), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_5103, signal_5102, signal_5101, signal_1837}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1823 ( .a ({signal_4260, signal_4259, signal_4258, signal_1556}), .b ({signal_4443, signal_4442, signal_4441, signal_1617}), .clk ( clk ), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({signal_5106, signal_5105, signal_5104, signal_1838}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1824 ( .a ({signal_3426, signal_3425, signal_3424, signal_1278}), .b ({signal_4668, signal_4667, signal_4666, signal_1692}), .clk ( clk ), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({signal_5109, signal_5108, signal_5107, signal_1839}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1825 ( .a ({signal_3306, signal_3305, signal_3304, signal_1238}), .b ({signal_4452, signal_4451, signal_4450, signal_1620}), .clk ( clk ), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({signal_5112, signal_5111, signal_5110, signal_1840}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1826 ( .a ({signal_3429, signal_3428, signal_3427, signal_1279}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({signal_5115, signal_5114, signal_5113, signal_1841}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1827 ( .a ({signal_3291, signal_3290, signal_3289, signal_1233}), .b ({signal_4677, signal_4676, signal_4675, signal_1695}), .clk ( clk ), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_5118, signal_5117, signal_5116, signal_1842}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1828 ( .a ({signal_4284, signal_4283, signal_4282, signal_1564}), .b ({signal_4461, signal_4460, signal_4459, signal_1623}), .clk ( clk ), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({signal_5121, signal_5120, signal_5119, signal_1843}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1829 ( .a ({signal_3450, signal_3449, signal_3448, signal_1286}), .b ({signal_4464, signal_4463, signal_4462, signal_1624}), .clk ( clk ), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({signal_5124, signal_5123, signal_5122, signal_1844}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1830 ( .a ({signal_4470, signal_4469, signal_4468, signal_1626}), .b ({signal_4473, signal_4472, signal_4471, signal_1627}), .clk ( clk ), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({signal_5127, signal_5126, signal_5125, signal_1845}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1831 ( .a ({signal_4368, signal_4367, signal_4366, signal_1592}), .b ({signal_4476, signal_4475, signal_4474, signal_1628}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({signal_5130, signal_5129, signal_5128, signal_1846}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1832 ( .a ({signal_4161, signal_4160, signal_4159, signal_1523}), .b ({signal_4494, signal_4493, signal_4492, signal_1634}), .clk ( clk ), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_5133, signal_5132, signal_5131, signal_1847}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1833 ( .a ({signal_3678, signal_3677, signal_3676, signal_1362}), .b ({signal_4497, signal_4496, signal_4495, signal_1635}), .clk ( clk ), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({signal_5136, signal_5135, signal_5134, signal_1848}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1842 ( .a ({signal_4926, signal_4925, signal_4924, signal_1778}), .b ({signal_5163, signal_5162, signal_5161, signal_1857}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1853 ( .a ({signal_4977, signal_4976, signal_4975, signal_1795}), .b ({signal_5196, signal_5195, signal_5194, signal_1868}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1859 ( .a ({signal_5007, signal_5006, signal_5005, signal_1805}), .b ({signal_5214, signal_5213, signal_5212, signal_1874}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1860 ( .a ({signal_5013, signal_5012, signal_5011, signal_1807}), .b ({signal_5217, signal_5216, signal_5215, signal_1875}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1861 ( .a ({signal_5028, signal_5027, signal_5026, signal_1812}), .b ({signal_5220, signal_5219, signal_5218, signal_1876}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1862 ( .a ({signal_5040, signal_5039, signal_5038, signal_1816}), .b ({signal_5223, signal_5222, signal_5221, signal_1877}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1863 ( .a ({signal_5043, signal_5042, signal_5041, signal_1817}), .b ({signal_5226, signal_5225, signal_5224, signal_1878}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1864 ( .a ({signal_5055, signal_5054, signal_5053, signal_1821}), .b ({signal_5229, signal_5228, signal_5227, signal_1879}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1865 ( .a ({signal_5058, signal_5057, signal_5056, signal_1822}), .b ({signal_5232, signal_5231, signal_5230, signal_1880}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1866 ( .a ({signal_5061, signal_5060, signal_5059, signal_1823}), .b ({signal_5235, signal_5234, signal_5233, signal_1881}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1867 ( .a ({signal_5064, signal_5063, signal_5062, signal_1824}), .b ({signal_5238, signal_5237, signal_5236, signal_1882}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1868 ( .a ({signal_5076, signal_5075, signal_5074, signal_1828}), .b ({signal_5241, signal_5240, signal_5239, signal_1883}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1869 ( .a ({signal_5079, signal_5078, signal_5077, signal_1829}), .b ({signal_5244, signal_5243, signal_5242, signal_1884}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1870 ( .a ({signal_5085, signal_5084, signal_5083, signal_1831}), .b ({signal_5247, signal_5246, signal_5245, signal_1885}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1871 ( .a ({signal_5088, signal_5087, signal_5086, signal_1832}), .b ({signal_5250, signal_5249, signal_5248, signal_1886}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1873 ( .a ({signal_5118, signal_5117, signal_5116, signal_1842}), .b ({signal_5256, signal_5255, signal_5254, signal_1888}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1874 ( .a ({signal_5124, signal_5123, signal_5122, signal_1844}), .b ({signal_5259, signal_5258, signal_5257, signal_1889}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1876 ( .a ({signal_4737, signal_4736, signal_4735, signal_1715}), .b ({signal_3387, signal_3386, signal_3385, signal_1265}), .clk ( clk ), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({signal_5265, signal_5264, signal_5263, signal_1891}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1877 ( .a ({signal_2466, signal_2465, signal_2464, signal_958}), .b ({signal_4740, signal_4739, signal_4738, signal_1716}), .clk ( clk ), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({signal_5268, signal_5267, signal_5266, signal_1892}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1878 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_4743, signal_4742, signal_4741, signal_1717}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({signal_5271, signal_5270, signal_5269, signal_1893}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1879 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_4746, signal_4745, signal_4744, signal_1718}), .clk ( clk ), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_5274, signal_5273, signal_5272, signal_1894}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1880 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_4896, signal_4895, signal_4894, signal_1768}), .clk ( clk ), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({signal_5277, signal_5276, signal_5275, signal_1895}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1881 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_4749, signal_4748, signal_4747, signal_1719}), .clk ( clk ), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({signal_5280, signal_5279, signal_5278, signal_1896}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1882 ( .a ({signal_4752, signal_4751, signal_4750, signal_1720}), .b ({signal_3591, signal_3590, signal_3589, signal_1333}), .clk ( clk ), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({signal_5283, signal_5282, signal_5281, signal_1897}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1883 ( .a ({signal_2613, signal_2612, signal_2611, signal_1007}), .b ({signal_4755, signal_4754, signal_4753, signal_1721}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({signal_5286, signal_5285, signal_5284, signal_1898}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1884 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({signal_4758, signal_4757, signal_4756, signal_1722}), .clk ( clk ), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_5289, signal_5288, signal_5287, signal_1899}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1885 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_4761, signal_4760, signal_4759, signal_1723}), .clk ( clk ), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({signal_5292, signal_5291, signal_5290, signal_1900}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1886 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_4899, signal_4898, signal_4897, signal_1769}), .clk ( clk ), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({signal_5295, signal_5294, signal_5293, signal_1901}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1887 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_4764, signal_4763, signal_4762, signal_1724}), .clk ( clk ), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({signal_5298, signal_5297, signal_5296, signal_1902}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1888 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_4770, signal_4769, signal_4768, signal_1726}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({signal_5301, signal_5300, signal_5299, signal_1903}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1889 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_4905, signal_4904, signal_4903, signal_1771}), .clk ( clk ), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_5304, signal_5303, signal_5302, signal_1904}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1890 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_4773, signal_4772, signal_4771, signal_1727}), .clk ( clk ), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({signal_5307, signal_5306, signal_5305, signal_1905}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1891 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_4776, signal_4775, signal_4774, signal_1728}), .clk ( clk ), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({signal_5310, signal_5309, signal_5308, signal_1906}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1892 ( .a ({signal_3027, signal_3026, signal_3025, signal_1145}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}), .clk ( clk ), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({signal_5313, signal_5312, signal_5311, signal_1907}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1894 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_4785, signal_4784, signal_4783, signal_1731}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({signal_5319, signal_5318, signal_5317, signal_1909}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1895 ( .a ({signal_2481, signal_2480, signal_2479, signal_963}), .b ({signal_4788, signal_4787, signal_4786, signal_1732}), .clk ( clk ), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_5322, signal_5321, signal_5320, signal_1910}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1896 ( .a ({signal_2877, signal_2876, signal_2875, signal_1095}), .b ({signal_4791, signal_4790, signal_4789, signal_1733}), .clk ( clk ), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({signal_5325, signal_5324, signal_5323, signal_1911}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1897 ( .a ({signal_2826, signal_2825, signal_2824, signal_1078}), .b ({signal_4794, signal_4793, signal_4792, signal_1734}), .clk ( clk ), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({signal_5328, signal_5327, signal_5326, signal_1912}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1898 ( .a ({signal_2811, signal_2810, signal_2809, signal_1073}), .b ({signal_4938, signal_4937, signal_4936, signal_1782}), .clk ( clk ), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({signal_5331, signal_5330, signal_5329, signal_1913}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1899 ( .a ({signal_3066, signal_3065, signal_3064, signal_1158}), .b ({signal_4797, signal_4796, signal_4795, signal_1735}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({signal_5334, signal_5333, signal_5332, signal_1914}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1900 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_4803, signal_4802, signal_4801, signal_1737}), .clk ( clk ), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_5337, signal_5336, signal_5335, signal_1915}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1901 ( .a ({signal_4806, signal_4805, signal_4804, signal_1738}), .b ({signal_4614, signal_4613, signal_4612, signal_1674}), .clk ( clk ), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({signal_5340, signal_5339, signal_5338, signal_1916}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1903 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_4809, signal_4808, signal_4807, signal_1739}), .clk ( clk ), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({signal_5346, signal_5345, signal_5344, signal_1918}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1905 ( .a ({signal_2877, signal_2876, signal_2875, signal_1095}), .b ({signal_4815, signal_4814, signal_4813, signal_1741}), .clk ( clk ), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({signal_5352, signal_5351, signal_5350, signal_1920}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1906 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_4818, signal_4817, signal_4816, signal_1742}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({signal_5355, signal_5354, signal_5353, signal_1921}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1907 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_4821, signal_4820, signal_4819, signal_1743}), .clk ( clk ), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_5358, signal_5357, signal_5356, signal_1922}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1908 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_4824, signal_4823, signal_4822, signal_1744}), .clk ( clk ), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({signal_5361, signal_5360, signal_5359, signal_1923}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1909 ( .a ({signal_2652, signal_2651, signal_2650, signal_1020}), .b ({signal_4938, signal_4937, signal_4936, signal_1782}), .clk ( clk ), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({signal_5364, signal_5363, signal_5362, signal_1924}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1910 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_4827, signal_4826, signal_4825, signal_1745}), .clk ( clk ), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({signal_5367, signal_5366, signal_5365, signal_1925}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1913 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_4830, signal_4829, signal_4828, signal_1746}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({signal_5376, signal_5375, signal_5374, signal_1928}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1914 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_4833, signal_4832, signal_4831, signal_1747}), .clk ( clk ), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_5379, signal_5378, signal_5377, signal_1929}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1915 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_4836, signal_4835, signal_4834, signal_1748}), .clk ( clk ), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({signal_5382, signal_5381, signal_5380, signal_1930}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1916 ( .a ({signal_3078, signal_3077, signal_3076, signal_1162}), .b ({signal_4767, signal_4766, signal_4765, signal_1725}), .clk ( clk ), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({signal_5385, signal_5384, signal_5383, signal_1931}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1917 ( .a ({signal_2805, signal_2804, signal_2803, signal_1071}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}), .clk ( clk ), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({signal_5388, signal_5387, signal_5386, signal_1932}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1919 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_4839, signal_4838, signal_4837, signal_1749}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({signal_5394, signal_5393, signal_5392, signal_1934}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1920 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_4842, signal_4841, signal_4840, signal_1750}), .clk ( clk ), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_5397, signal_5396, signal_5395, signal_1935}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1923 ( .a ({signal_2835, signal_2834, signal_2833, signal_1081}), .b ({signal_4845, signal_4844, signal_4843, signal_1751}), .clk ( clk ), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({signal_5406, signal_5405, signal_5404, signal_1938}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1927 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_4854, signal_4853, signal_4852, signal_1754}), .clk ( clk ), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({signal_5418, signal_5417, signal_5416, signal_1942}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1932 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_4872, signal_4871, signal_4870, signal_1760}), .clk ( clk ), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({signal_5433, signal_5432, signal_5431, signal_1947}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1944 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_4884, signal_4883, signal_4882, signal_1764}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({signal_5469, signal_5468, signal_5467, signal_1959}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1948 ( .a ({signal_5268, signal_5267, signal_5266, signal_1892}), .b ({signal_5481, signal_5480, signal_5479, signal_1963}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1949 ( .a ({signal_5271, signal_5270, signal_5269, signal_1893}), .b ({signal_5484, signal_5483, signal_5482, signal_1964}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1950 ( .a ({signal_5277, signal_5276, signal_5275, signal_1895}), .b ({signal_5487, signal_5486, signal_5485, signal_1965}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1951 ( .a ({signal_5283, signal_5282, signal_5281, signal_1897}), .b ({signal_5490, signal_5489, signal_5488, signal_1966}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1952 ( .a ({signal_5286, signal_5285, signal_5284, signal_1898}), .b ({signal_5493, signal_5492, signal_5491, signal_1967}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1953 ( .a ({signal_5292, signal_5291, signal_5290, signal_1900}), .b ({signal_5496, signal_5495, signal_5494, signal_1968}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1954 ( .a ({signal_5295, signal_5294, signal_5293, signal_1901}), .b ({signal_5499, signal_5498, signal_5497, signal_1969}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1955 ( .a ({signal_5298, signal_5297, signal_5296, signal_1902}), .b ({signal_5502, signal_5501, signal_5500, signal_1970}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1956 ( .a ({signal_5301, signal_5300, signal_5299, signal_1903}), .b ({signal_5505, signal_5504, signal_5503, signal_1971}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1957 ( .a ({signal_5304, signal_5303, signal_5302, signal_1904}), .b ({signal_5508, signal_5507, signal_5506, signal_1972}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1958 ( .a ({signal_5307, signal_5306, signal_5305, signal_1905}), .b ({signal_5511, signal_5510, signal_5509, signal_1973}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1959 ( .a ({signal_5310, signal_5309, signal_5308, signal_1906}), .b ({signal_5514, signal_5513, signal_5512, signal_1974}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1960 ( .a ({signal_5313, signal_5312, signal_5311, signal_1907}), .b ({signal_5517, signal_5516, signal_5515, signal_1975}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1962 ( .a ({signal_5319, signal_5318, signal_5317, signal_1909}), .b ({signal_5523, signal_5522, signal_5521, signal_1977}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1963 ( .a ({signal_5322, signal_5321, signal_5320, signal_1910}), .b ({signal_5526, signal_5525, signal_5524, signal_1978}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1964 ( .a ({signal_5325, signal_5324, signal_5323, signal_1911}), .b ({signal_5529, signal_5528, signal_5527, signal_1979}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1965 ( .a ({signal_5328, signal_5327, signal_5326, signal_1912}), .b ({signal_5532, signal_5531, signal_5530, signal_1980}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1966 ( .a ({signal_5331, signal_5330, signal_5329, signal_1913}), .b ({signal_5535, signal_5534, signal_5533, signal_1981}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1967 ( .a ({signal_5334, signal_5333, signal_5332, signal_1914}), .b ({signal_5538, signal_5537, signal_5536, signal_1982}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1968 ( .a ({signal_5337, signal_5336, signal_5335, signal_1915}), .b ({signal_5541, signal_5540, signal_5539, signal_1983}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1970 ( .a ({signal_5346, signal_5345, signal_5344, signal_1918}), .b ({signal_5547, signal_5546, signal_5545, signal_1985}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1972 ( .a ({signal_5352, signal_5351, signal_5350, signal_1920}), .b ({signal_5553, signal_5552, signal_5551, signal_1987}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1973 ( .a ({signal_5355, signal_5354, signal_5353, signal_1921}), .b ({signal_5556, signal_5555, signal_5554, signal_1988}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1974 ( .a ({signal_5358, signal_5357, signal_5356, signal_1922}), .b ({signal_5559, signal_5558, signal_5557, signal_1989}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1975 ( .a ({signal_5361, signal_5360, signal_5359, signal_1923}), .b ({signal_5562, signal_5561, signal_5560, signal_1990}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1976 ( .a ({signal_5364, signal_5363, signal_5362, signal_1924}), .b ({signal_5565, signal_5564, signal_5563, signal_1991}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1977 ( .a ({signal_5367, signal_5366, signal_5365, signal_1925}), .b ({signal_5568, signal_5567, signal_5566, signal_1992}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1979 ( .a ({signal_5376, signal_5375, signal_5374, signal_1928}), .b ({signal_5574, signal_5573, signal_5572, signal_1994}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1980 ( .a ({signal_5379, signal_5378, signal_5377, signal_1929}), .b ({signal_5577, signal_5576, signal_5575, signal_1995}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1981 ( .a ({signal_5382, signal_5381, signal_5380, signal_1930}), .b ({signal_5580, signal_5579, signal_5578, signal_1996}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1982 ( .a ({signal_5385, signal_5384, signal_5383, signal_1931}), .b ({signal_5583, signal_5582, signal_5581, signal_1997}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1983 ( .a ({signal_5388, signal_5387, signal_5386, signal_1932}), .b ({signal_5586, signal_5585, signal_5584, signal_1998}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1984 ( .a ({signal_5394, signal_5393, signal_5392, signal_1934}), .b ({signal_5589, signal_5588, signal_5587, signal_1999}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1985 ( .a ({signal_5397, signal_5396, signal_5395, signal_1935}), .b ({signal_5592, signal_5591, signal_5590, signal_2000}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1988 ( .a ({signal_5406, signal_5405, signal_5404, signal_1938}), .b ({signal_5601, signal_5600, signal_5599, signal_2003}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1990 ( .a ({signal_5418, signal_5417, signal_5416, signal_1942}), .b ({signal_5607, signal_5606, signal_5605, signal_2005}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1991 ( .a ({signal_5433, signal_5432, signal_5431, signal_1947}), .b ({signal_5610, signal_5609, signal_5608, signal_2006}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1996 ( .a ({signal_5469, signal_5468, signal_5467, signal_1959}), .b ({signal_5625, signal_5624, signal_5623, signal_2011}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2000 ( .a ({signal_5181, signal_5180, signal_5179, signal_1863}), .b ({signal_4374, signal_4373, signal_4372, signal_1594}), .clk ( clk ), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_5637, signal_5636, signal_5635, signal_2015}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2001 ( .a ({signal_5148, signal_5147, signal_5146, signal_1852}), .b ({signal_4287, signal_4286, signal_4285, signal_1565}), .clk ( clk ), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({signal_5640, signal_5639, signal_5638, signal_2016}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2003 ( .a ({signal_5157, signal_5156, signal_5155, signal_1855}), .b ({signal_5160, signal_5159, signal_5158, signal_1856}), .clk ( clk ), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({signal_5646, signal_5645, signal_5644, signal_2018}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2004 ( .a ({signal_3504, signal_3503, signal_3502, signal_1304}), .b ({signal_5166, signal_5165, signal_5164, signal_1858}), .clk ( clk ), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({signal_5649, signal_5648, signal_5647, signal_2019}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2005 ( .a ({signal_2778, signal_2777, signal_2776, signal_1062}), .b ({signal_5169, signal_5168, signal_5167, signal_1859}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({signal_5652, signal_5651, signal_5650, signal_2020}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2006 ( .a ({signal_3342, signal_3341, signal_3340, signal_1250}), .b ({signal_5172, signal_5171, signal_5170, signal_1860}), .clk ( clk ), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_5655, signal_5654, signal_5653, signal_2021}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2008 ( .a ({signal_3573, signal_3572, signal_3571, signal_1327}), .b ({signal_5184, signal_5183, signal_5182, signal_1864}), .clk ( clk ), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({signal_5661, signal_5660, signal_5659, signal_2023}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2011 ( .a ({signal_2778, signal_2777, signal_2776, signal_1062}), .b ({signal_5187, signal_5186, signal_5185, signal_1865}), .clk ( clk ), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({signal_5670, signal_5669, signal_5668, signal_2026}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2012 ( .a ({signal_4419, signal_4418, signal_4417, signal_1609}), .b ({signal_5193, signal_5192, signal_5191, signal_1867}), .clk ( clk ), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({signal_5673, signal_5672, signal_5671, signal_2027}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2014 ( .a ({signal_5199, signal_5198, signal_5197, signal_1869}), .b ({signal_4656, signal_4655, signal_4654, signal_1688}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({signal_5679, signal_5678, signal_5677, signal_2029}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2015 ( .a ({signal_4413, signal_4412, signal_4411, signal_1607}), .b ({signal_5205, signal_5204, signal_5203, signal_1871}), .clk ( clk ), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_5682, signal_5681, signal_5680, signal_2030}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2048 ( .a ({signal_5649, signal_5648, signal_5647, signal_2019}), .b ({signal_5781, signal_5780, signal_5779, signal_2063}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2052 ( .a ({signal_5670, signal_5669, signal_5668, signal_2026}), .b ({signal_5793, signal_5792, signal_5791, signal_2067}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1819 ( .a ({signal_4242, signal_4241, signal_4240, signal_1550}), .b ({signal_4653, signal_4652, signal_4651, signal_1687}), .clk ( clk ), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({signal_5094, signal_5093, signal_5092, signal_1834}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1834 ( .a ({signal_4290, signal_4289, signal_4288, signal_1566}), .b ({signal_4722, signal_4721, signal_4720, signal_1710}), .clk ( clk ), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({signal_5139, signal_5138, signal_5137, signal_1849}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1872 ( .a ({signal_5094, signal_5093, signal_5092, signal_1834}), .b ({signal_5253, signal_5252, signal_5251, signal_1887}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1875 ( .a ({signal_5139, signal_5138, signal_5137, signal_1849}), .b ({signal_5262, signal_5261, signal_5260, signal_1890}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1893 ( .a ({signal_2574, signal_2573, signal_2572, signal_994}), .b ({signal_4782, signal_4781, signal_4780, signal_1730}), .clk ( clk ), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({signal_5316, signal_5315, signal_5314, signal_1908}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1902 ( .a ({signal_4893, signal_4892, signal_4891, signal_1767}), .b ({signal_4950, signal_4949, signal_4948, signal_1786}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({signal_5343, signal_5342, signal_5341, signal_1917}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1904 ( .a ({signal_2574, signal_2573, signal_2572, signal_994}), .b ({signal_4812, signal_4811, signal_4810, signal_1740}), .clk ( clk ), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_5349, signal_5348, signal_5347, signal_1919}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1911 ( .a ({signal_4962, signal_4961, signal_4960, signal_1790}), .b ({signal_4404, signal_4403, signal_4402, signal_1604}), .clk ( clk ), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({signal_5370, signal_5369, signal_5368, signal_1926}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1912 ( .a ({signal_3462, signal_3461, signal_3460, signal_1290}), .b ({signal_4968, signal_4967, signal_4966, signal_1792}), .clk ( clk ), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({signal_5373, signal_5372, signal_5371, signal_1927}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1918 ( .a ({signal_3654, signal_3653, signal_3652, signal_1354}), .b ({signal_5004, signal_5003, signal_5002, signal_1804}), .clk ( clk ), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({signal_5391, signal_5390, signal_5389, signal_1933}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1921 ( .a ({signal_3294, signal_3293, signal_3292, signal_1234}), .b ({signal_5010, signal_5009, signal_5008, signal_1806}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({signal_5400, signal_5399, signal_5398, signal_1936}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1922 ( .a ({signal_5016, signal_5015, signal_5014, signal_1808}), .b ({signal_5019, signal_5018, signal_5017, signal_1809}), .clk ( clk ), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_5403, signal_5402, signal_5401, signal_1937}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1924 ( .a ({signal_2523, signal_2522, signal_2521, signal_977}), .b ({signal_4848, signal_4847, signal_4846, signal_1752}), .clk ( clk ), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({signal_5409, signal_5408, signal_5407, signal_1939}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1925 ( .a ({signal_4320, signal_4319, signal_4318, signal_1576}), .b ({signal_5037, signal_5036, signal_5035, signal_1815}), .clk ( clk ), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({signal_5412, signal_5411, signal_5410, signal_1940}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1926 ( .a ({signal_4338, signal_4337, signal_4336, signal_1582}), .b ({signal_4851, signal_4850, signal_4849, signal_1753}), .clk ( clk ), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({signal_5415, signal_5414, signal_5413, signal_1941}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1928 ( .a ({signal_3531, signal_3530, signal_3529, signal_1313}), .b ({signal_5049, signal_5048, signal_5047, signal_1819}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({signal_5421, signal_5420, signal_5419, signal_1943}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1929 ( .a ({signal_4959, signal_4958, signal_4957, signal_1789}), .b ({signal_4488, signal_4487, signal_4486, signal_1632}), .clk ( clk ), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_5424, signal_5423, signal_5422, signal_1944}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1930 ( .a ({signal_4860, signal_4859, signal_4858, signal_1756}), .b ({signal_4863, signal_4862, signal_4861, signal_1757}), .clk ( clk ), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({signal_5427, signal_5426, signal_5425, signal_1945}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1931 ( .a ({signal_4383, signal_4382, signal_4381, signal_1597}), .b ({signal_4869, signal_4868, signal_4867, signal_1759}), .clk ( clk ), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({signal_5430, signal_5429, signal_5428, signal_1946}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1933 ( .a ({signal_3597, signal_3596, signal_3595, signal_1335}), .b ({signal_5073, signal_5072, signal_5071, signal_1827}), .clk ( clk ), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({signal_5436, signal_5435, signal_5434, signal_1948}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1934 ( .a ({signal_4377, signal_4376, signal_4375, signal_1595}), .b ({signal_5091, signal_5090, signal_5089, signal_1833}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({signal_5439, signal_5438, signal_5437, signal_1949}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1935 ( .a ({signal_4245, signal_4244, signal_4243, signal_1551}), .b ({signal_5097, signal_5096, signal_5095, signal_1835}), .clk ( clk ), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_5442, signal_5441, signal_5440, signal_1950}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1936 ( .a ({signal_4875, signal_4874, signal_4873, signal_1761}), .b ({signal_5100, signal_5099, signal_5098, signal_1836}), .clk ( clk ), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({signal_5445, signal_5444, signal_5443, signal_1951}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1937 ( .a ({signal_4431, signal_4430, signal_4429, signal_1613}), .b ({signal_4857, signal_4856, signal_4855, signal_1755}), .clk ( clk ), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({signal_5448, signal_5447, signal_5446, signal_1952}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1938 ( .a ({signal_4662, signal_4661, signal_4660, signal_1690}), .b ({signal_5103, signal_5102, signal_5101, signal_1837}), .clk ( clk ), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({signal_5451, signal_5450, signal_5449, signal_1953}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1939 ( .a ({signal_4257, signal_4256, signal_4255, signal_1555}), .b ({signal_5106, signal_5105, signal_5104, signal_1838}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({signal_5454, signal_5453, signal_5452, signal_1954}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1940 ( .a ({signal_2775, signal_2774, signal_2773, signal_1061}), .b ({signal_5112, signal_5111, signal_5110, signal_1840}), .clk ( clk ), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_5457, signal_5456, signal_5455, signal_1955}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1941 ( .a ({signal_4278, signal_4277, signal_4276, signal_1562}), .b ({signal_4881, signal_4880, signal_4879, signal_1763}), .clk ( clk ), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({signal_5460, signal_5459, signal_5458, signal_1956}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1942 ( .a ({signal_4674, signal_4673, signal_4672, signal_1694}), .b ({signal_5115, signal_5114, signal_5113, signal_1841}), .clk ( clk ), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({signal_5463, signal_5462, signal_5461, signal_1957}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1943 ( .a ({signal_5001, signal_5000, signal_4999, signal_1803}), .b ({signal_4500, signal_4499, signal_4498, signal_1636}), .clk ( clk ), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({signal_5466, signal_5465, signal_5464, signal_1958}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1945 ( .a ({signal_5067, signal_5066, signal_5065, signal_1825}), .b ({signal_5130, signal_5129, signal_5128, signal_1846}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({signal_5472, signal_5471, signal_5470, signal_1960}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1946 ( .a ({signal_4296, signal_4295, signal_4294, signal_1568}), .b ({signal_4887, signal_4886, signal_4885, signal_1765}), .clk ( clk ), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_5475, signal_5474, signal_5473, signal_1961}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1947 ( .a ({signal_4980, signal_4979, signal_4978, signal_1796}), .b ({signal_5133, signal_5132, signal_5131, signal_1847}), .clk ( clk ), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({signal_5478, signal_5477, signal_5476, signal_1962}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1961 ( .a ({signal_5316, signal_5315, signal_5314, signal_1908}), .b ({signal_5520, signal_5519, signal_5518, signal_1976}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1969 ( .a ({signal_5343, signal_5342, signal_5341, signal_1917}), .b ({signal_5544, signal_5543, signal_5542, signal_1984}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1971 ( .a ({signal_5349, signal_5348, signal_5347, signal_1919}), .b ({signal_5550, signal_5549, signal_5548, signal_1986}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1978 ( .a ({signal_5373, signal_5372, signal_5371, signal_1927}), .b ({signal_5571, signal_5570, signal_5569, signal_1993}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1986 ( .a ({signal_5400, signal_5399, signal_5398, signal_1936}), .b ({signal_5595, signal_5594, signal_5593, signal_2001}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1987 ( .a ({signal_5403, signal_5402, signal_5401, signal_1937}), .b ({signal_5598, signal_5597, signal_5596, signal_2002}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1989 ( .a ({signal_5409, signal_5408, signal_5407, signal_1939}), .b ({signal_5604, signal_5603, signal_5602, signal_2004}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1992 ( .a ({signal_5439, signal_5438, signal_5437, signal_1949}), .b ({signal_5613, signal_5612, signal_5611, signal_2007}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1993 ( .a ({signal_5445, signal_5444, signal_5443, signal_1951}), .b ({signal_5616, signal_5615, signal_5614, signal_2008}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1994 ( .a ({signal_5463, signal_5462, signal_5461, signal_1957}), .b ({signal_5619, signal_5618, signal_5617, signal_2009}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1995 ( .a ({signal_5466, signal_5465, signal_5464, signal_1958}), .b ({signal_5622, signal_5621, signal_5620, signal_2010}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1997 ( .a ({signal_5472, signal_5471, signal_5470, signal_1960}), .b ({signal_5628, signal_5627, signal_5626, signal_2012}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_1998 ( .a ({signal_5478, signal_5477, signal_5476, signal_1962}), .b ({signal_5631, signal_5630, signal_5629, signal_2013}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_1999 ( .a ({signal_5163, signal_5162, signal_5161, signal_1857}), .b ({signal_3675, signal_3674, signal_3673, signal_1361}), .clk ( clk ), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({signal_5634, signal_5633, signal_5632, signal_2014}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2002 ( .a ({signal_5151, signal_5150, signal_5149, signal_1853}), .b ({signal_4914, signal_4913, signal_4912, signal_1774}), .clk ( clk ), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({signal_5643, signal_5642, signal_5641, signal_2017}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2007 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_5274, signal_5273, signal_5272, signal_1894}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({signal_5658, signal_5657, signal_5656, signal_2022}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2009 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_5280, signal_5279, signal_5278, signal_1896}), .clk ( clk ), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_5664, signal_5663, signal_5662, signal_2024}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2010 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_5289, signal_5288, signal_5287, signal_1899}), .clk ( clk ), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({signal_5667, signal_5666, signal_5665, signal_2025}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2013 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_5196, signal_5195, signal_5194, signal_1868}), .clk ( clk ), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({signal_5676, signal_5675, signal_5674, signal_2028}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2016 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_5214, signal_5213, signal_5212, signal_1874}), .clk ( clk ), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({signal_5685, signal_5684, signal_5683, signal_2031}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2017 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_5217, signal_5216, signal_5215, signal_1875}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({signal_5688, signal_5687, signal_5686, signal_2032}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2018 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_5220, signal_5219, signal_5218, signal_1876}), .clk ( clk ), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_5691, signal_5690, signal_5689, signal_2033}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2019 ( .a ({signal_5154, signal_5153, signal_5152, signal_1854}), .b ({signal_5031, signal_5030, signal_5029, signal_1813}), .clk ( clk ), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({signal_5694, signal_5693, signal_5692, signal_2034}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2020 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_5223, signal_5222, signal_5221, signal_1877}), .clk ( clk ), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({signal_5697, signal_5696, signal_5695, signal_2035}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2021 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_5226, signal_5225, signal_5224, signal_1878}), .clk ( clk ), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({signal_5700, signal_5699, signal_5698, signal_2036}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2022 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_5229, signal_5228, signal_5227, signal_1879}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({signal_5703, signal_5702, signal_5701, signal_2037}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2023 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_5232, signal_5231, signal_5230, signal_1880}), .clk ( clk ), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_5706, signal_5705, signal_5704, signal_2038}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2024 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_5235, signal_5234, signal_5233, signal_1881}), .clk ( clk ), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({signal_5709, signal_5708, signal_5707, signal_2039}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2025 ( .a ({signal_5178, signal_5177, signal_5176, signal_1862}), .b ({signal_5238, signal_5237, signal_5236, signal_1882}), .clk ( clk ), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({signal_5712, signal_5711, signal_5710, signal_2040}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2026 ( .a ({signal_5070, signal_5069, signal_5068, signal_1826}), .b ({signal_5340, signal_5339, signal_5338, signal_1916}), .clk ( clk ), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({signal_5715, signal_5714, signal_5713, signal_2041}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2028 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_5241, signal_5240, signal_5239, signal_1883}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({signal_5721, signal_5720, signal_5719, signal_2043}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2029 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_5244, signal_5243, signal_5242, signal_1884}), .clk ( clk ), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_5724, signal_5723, signal_5722, signal_2044}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2030 ( .a ({signal_5190, signal_5189, signal_5188, signal_1866}), .b ({signal_5082, signal_5081, signal_5080, signal_1830}), .clk ( clk ), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({signal_5727, signal_5726, signal_5725, signal_2045}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2031 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_5250, signal_5249, signal_5248, signal_1886}), .clk ( clk ), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({signal_5730, signal_5729, signal_5728, signal_2046}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2033 ( .a ({signal_5211, signal_5210, signal_5209, signal_1873}), .b ({signal_5109, signal_5108, signal_5107, signal_1839}), .clk ( clk ), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({signal_5736, signal_5735, signal_5734, signal_2048}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2034 ( .a ({signal_5145, signal_5144, signal_5143, signal_1851}), .b ({signal_5046, signal_5045, signal_5044, signal_1818}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({signal_5739, signal_5738, signal_5737, signal_2049}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2035 ( .a ({signal_2832, signal_2831, signal_2830, signal_1080}), .b ({signal_5256, signal_5255, signal_5254, signal_1888}), .clk ( clk ), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_5742, signal_5741, signal_5740, signal_2050}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2036 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_5259, signal_5258, signal_5257, signal_1889}), .clk ( clk ), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({signal_5745, signal_5744, signal_5743, signal_2051}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2046 ( .a ({signal_5634, signal_5633, signal_5632, signal_2014}), .b ({signal_5775, signal_5774, signal_5773, signal_2061}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2047 ( .a ({signal_5643, signal_5642, signal_5641, signal_2017}), .b ({signal_5778, signal_5777, signal_5776, signal_2062}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2049 ( .a ({signal_5658, signal_5657, signal_5656, signal_2022}), .b ({signal_5784, signal_5783, signal_5782, signal_2064}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2050 ( .a ({signal_5664, signal_5663, signal_5662, signal_2024}), .b ({signal_5787, signal_5786, signal_5785, signal_2065}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2051 ( .a ({signal_5667, signal_5666, signal_5665, signal_2025}), .b ({signal_5790, signal_5789, signal_5788, signal_2066}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2053 ( .a ({signal_5676, signal_5675, signal_5674, signal_2028}), .b ({signal_5796, signal_5795, signal_5794, signal_2068}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2054 ( .a ({signal_5685, signal_5684, signal_5683, signal_2031}), .b ({signal_5799, signal_5798, signal_5797, signal_2069}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2055 ( .a ({signal_5688, signal_5687, signal_5686, signal_2032}), .b ({signal_5802, signal_5801, signal_5800, signal_2070}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2056 ( .a ({signal_5691, signal_5690, signal_5689, signal_2033}), .b ({signal_5805, signal_5804, signal_5803, signal_2071}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2057 ( .a ({signal_5694, signal_5693, signal_5692, signal_2034}), .b ({signal_5808, signal_5807, signal_5806, signal_2072}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2058 ( .a ({signal_5697, signal_5696, signal_5695, signal_2035}), .b ({signal_5811, signal_5810, signal_5809, signal_2073}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2059 ( .a ({signal_5700, signal_5699, signal_5698, signal_2036}), .b ({signal_5814, signal_5813, signal_5812, signal_2074}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2060 ( .a ({signal_5703, signal_5702, signal_5701, signal_2037}), .b ({signal_5817, signal_5816, signal_5815, signal_2075}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2061 ( .a ({signal_5706, signal_5705, signal_5704, signal_2038}), .b ({signal_5820, signal_5819, signal_5818, signal_2076}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2062 ( .a ({signal_5709, signal_5708, signal_5707, signal_2039}), .b ({signal_5823, signal_5822, signal_5821, signal_2077}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2063 ( .a ({signal_5715, signal_5714, signal_5713, signal_2041}), .b ({signal_5826, signal_5825, signal_5824, signal_2078}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2065 ( .a ({signal_5721, signal_5720, signal_5719, signal_2043}), .b ({signal_5832, signal_5831, signal_5830, signal_2080}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2066 ( .a ({signal_5724, signal_5723, signal_5722, signal_2044}), .b ({signal_5835, signal_5834, signal_5833, signal_2081}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2067 ( .a ({signal_5730, signal_5729, signal_5728, signal_2046}), .b ({signal_5838, signal_5837, signal_5836, signal_2082}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2069 ( .a ({signal_5736, signal_5735, signal_5734, signal_2048}), .b ({signal_5844, signal_5843, signal_5842, signal_2084}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2070 ( .a ({signal_5742, signal_5741, signal_5740, signal_2050}), .b ({signal_5847, signal_5846, signal_5845, signal_2085}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2071 ( .a ({signal_5745, signal_5744, signal_5743, signal_2051}), .b ({signal_5850, signal_5849, signal_5848, signal_2086}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2074 ( .a ({signal_5523, signal_5522, signal_5521, signal_1977}), .b ({signal_3687, signal_3686, signal_3685, signal_1365}), .clk ( clk ), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({signal_5859, signal_5858, signal_5857, signal_2089}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2075 ( .a ({signal_4305, signal_4304, signal_4303, signal_1571}), .b ({signal_5484, signal_5483, signal_5482, signal_1964}), .clk ( clk ), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({signal_5862, signal_5861, signal_5860, signal_2090}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2076 ( .a ({signal_3318, signal_3317, signal_3316, signal_1242}), .b ({signal_5637, signal_5636, signal_5635, signal_2015}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({signal_5865, signal_5864, signal_5863, signal_2091}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2077 ( .a ({signal_4212, signal_4211, signal_4210, signal_1540}), .b ({signal_5499, signal_5498, signal_5497, signal_1969}), .clk ( clk ), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_5868, signal_5867, signal_5866, signal_2092}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2078 ( .a ({signal_5481, signal_5480, signal_5479, signal_1963}), .b ({signal_5208, signal_5207, signal_5206, signal_1872}), .clk ( clk ), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({signal_5871, signal_5870, signal_5869, signal_2093}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2079 ( .a ({signal_5511, signal_5510, signal_5509, signal_1973}), .b ({signal_5514, signal_5513, signal_5512, signal_1974}), .clk ( clk ), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({signal_5874, signal_5873, signal_5872, signal_2094}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2080 ( .a ({signal_3480, signal_3479, signal_3478, signal_1296}), .b ({signal_5646, signal_5645, signal_5644, signal_2018}), .clk ( clk ), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({signal_5877, signal_5876, signal_5875, signal_2095}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2081 ( .a ({signal_3516, signal_3515, signal_3514, signal_1308}), .b ({signal_5652, signal_5651, signal_5650, signal_2020}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({signal_5880, signal_5879, signal_5878, signal_2096}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2082 ( .a ({signal_3345, signal_3344, signal_3343, signal_1251}), .b ({signal_5655, signal_5654, signal_5653, signal_2021}), .clk ( clk ), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_5883, signal_5882, signal_5881, signal_2097}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2083 ( .a ({signal_4341, signal_4340, signal_4339, signal_1583}), .b ({signal_5535, signal_5534, signal_5533, signal_1981}), .clk ( clk ), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({signal_5886, signal_5885, signal_5884, signal_2098}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2085 ( .a ({signal_3570, signal_3569, signal_3568, signal_1326}), .b ({signal_5547, signal_5546, signal_5545, signal_1985}), .clk ( clk ), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({signal_5892, signal_5891, signal_5890, signal_2100}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2086 ( .a ({signal_3375, signal_3374, signal_3373, signal_1261}), .b ({signal_5661, signal_5660, signal_5659, signal_2023}), .clk ( clk ), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({signal_5895, signal_5894, signal_5893, signal_2101}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2087 ( .a ({signal_5265, signal_5264, signal_5263, signal_1891}), .b ({signal_5559, signal_5558, signal_5557, signal_1989}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({signal_5898, signal_5897, signal_5896, signal_2102}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2088 ( .a ({signal_5562, signal_5561, signal_5560, signal_1990}), .b ({signal_5565, signal_5564, signal_5563, signal_1991}), .clk ( clk ), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_5901, signal_5900, signal_5899, signal_2103}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2089 ( .a ({signal_4392, signal_4391, signal_4390, signal_1600}), .b ({signal_5568, signal_5567, signal_5566, signal_1992}), .clk ( clk ), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({signal_5904, signal_5903, signal_5902, signal_2104}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2091 ( .a ({signal_5673, signal_5672, signal_5671, signal_2027}), .b ({signal_5247, signal_5246, signal_5245, signal_1885}), .clk ( clk ), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({signal_5910, signal_5909, signal_5908, signal_2106}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2092 ( .a ({signal_3405, signal_3404, signal_3403, signal_1271}), .b ({signal_5574, signal_5573, signal_5572, signal_1994}), .clk ( clk ), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({signal_5913, signal_5912, signal_5911, signal_2107}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2093 ( .a ({signal_5202, signal_5201, signal_5200, signal_1870}), .b ({signal_5577, signal_5576, signal_5575, signal_1995}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({signal_5916, signal_5915, signal_5914, signal_2108}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2094 ( .a ({signal_4998, signal_4997, signal_4996, signal_1802}), .b ({signal_5580, signal_5579, signal_5578, signal_1996}), .clk ( clk ), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_5919, signal_5918, signal_5917, signal_2109}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2095 ( .a ({signal_5505, signal_5504, signal_5503, signal_1971}), .b ({signal_5583, signal_5582, signal_5581, signal_1997}), .clk ( clk ), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({signal_5922, signal_5921, signal_5920, signal_2110}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2096 ( .a ({signal_4860, signal_4859, signal_4858, signal_1756}), .b ({signal_5586, signal_5585, signal_5584, signal_1998}), .clk ( clk ), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({signal_5925, signal_5924, signal_5923, signal_2111}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2097 ( .a ({signal_5508, signal_5507, signal_5506, signal_1972}), .b ({signal_4488, signal_4487, signal_4486, signal_1632}), .clk ( clk ), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({signal_5928, signal_5927, signal_5926, signal_2112}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2099 ( .a ({signal_4686, signal_4685, signal_4684, signal_1698}), .b ({signal_5592, signal_5591, signal_5590, signal_2000}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({signal_5934, signal_5933, signal_5932, signal_2114}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2101 ( .a ({signal_5517, signal_5516, signal_5515, signal_1975}), .b ({signal_5601, signal_5600, signal_5599, signal_2003}), .clk ( clk ), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_5940, signal_5939, signal_5938, signal_2116}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2104 ( .a ({signal_3528, signal_3527, signal_3526, signal_1312}), .b ({signal_5607, signal_5606, signal_5605, signal_2005}), .clk ( clk ), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({signal_5949, signal_5948, signal_5947, signal_2119}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2110 ( .a ({signal_5679, signal_5678, signal_5677, signal_2029}), .b ({signal_5136, signal_5135, signal_5134, signal_1848}), .clk ( clk ), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({signal_5967, signal_5966, signal_5965, signal_2125}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2124 ( .a ({signal_5859, signal_5858, signal_5857, signal_2089}), .b ({signal_6009, signal_6008, signal_6007, signal_2139}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2125 ( .a ({signal_5865, signal_5864, signal_5863, signal_2091}), .b ({signal_6012, signal_6011, signal_6010, signal_2140}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2126 ( .a ({signal_5868, signal_5867, signal_5866, signal_2092}), .b ({signal_6015, signal_6014, signal_6013, signal_2141}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2127 ( .a ({signal_5880, signal_5879, signal_5878, signal_2096}), .b ({signal_6018, signal_6017, signal_6016, signal_2142}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2128 ( .a ({signal_5883, signal_5882, signal_5881, signal_2097}), .b ({signal_6021, signal_6020, signal_6019, signal_2143}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2130 ( .a ({signal_5895, signal_5894, signal_5893, signal_2101}), .b ({signal_6027, signal_6026, signal_6025, signal_2145}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2133 ( .a ({signal_5949, signal_5948, signal_5947, signal_2119}), .b ({signal_6036, signal_6035, signal_6034, signal_2148}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2135 ( .a ({signal_5967, signal_5966, signal_5965, signal_2125}), .b ({signal_6042, signal_6041, signal_6040, signal_2150}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2144 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_5781, signal_5780, signal_5779, signal_2063}), .clk ( clk ), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({signal_6069, signal_6068, signal_6067, signal_2159}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2148 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_5793, signal_5792, signal_5791, signal_2067}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({signal_6081, signal_6080, signal_6079, signal_2163}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2185 ( .a ({signal_6069, signal_6068, signal_6067, signal_2159}), .b ({signal_6192, signal_6191, signal_6190, signal_2200}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2186 ( .a ({signal_6081, signal_6080, signal_6079, signal_2163}), .b ({signal_6195, signal_6194, signal_6193, signal_2201}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2027 ( .a ({signal_4212, signal_4211, signal_4210, signal_1540}), .b ({signal_5370, signal_5369, signal_5368, signal_1926}), .clk ( clk ), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_5718, signal_5717, signal_5716, signal_2042}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2032 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_5253, signal_5252, signal_5251, signal_1887}), .clk ( clk ), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({signal_5733, signal_5732, signal_5731, signal_2047}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2037 ( .a ({signal_3336, signal_3335, signal_3334, signal_1248}), .b ({signal_5412, signal_5411, signal_5410, signal_1940}), .clk ( clk ), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({signal_5748, signal_5747, signal_5746, signal_2052}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2038 ( .a ({signal_3534, signal_3533, signal_3532, signal_1314}), .b ({signal_5421, signal_5420, signal_5419, signal_1943}), .clk ( clk ), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({signal_5751, signal_5750, signal_5749, signal_2053}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2039 ( .a ({signal_4203, signal_4202, signal_4201, signal_1537}), .b ({signal_5430, signal_5429, signal_5428, signal_1946}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({signal_5754, signal_5753, signal_5752, signal_2054}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2040 ( .a ({signal_3600, signal_3599, signal_3598, signal_1336}), .b ({signal_5436, signal_5435, signal_5434, signal_1948}), .clk ( clk ), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_5757, signal_5756, signal_5755, signal_2055}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2041 ( .a ({signal_4248, signal_4247, signal_4246, signal_1552}), .b ({signal_5442, signal_5441, signal_5440, signal_1950}), .clk ( clk ), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({signal_5760, signal_5759, signal_5758, signal_2056}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2042 ( .a ({signal_4446, signal_4445, signal_4444, signal_1618}), .b ({signal_5454, signal_5453, signal_5452, signal_1954}), .clk ( clk ), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({signal_5763, signal_5762, signal_5761, signal_2057}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2043 ( .a ({signal_4272, signal_4271, signal_4270, signal_1560}), .b ({signal_5457, signal_5456, signal_5455, signal_1955}), .clk ( clk ), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({signal_5766, signal_5765, signal_5764, signal_2058}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2044 ( .a ({signal_4458, signal_4457, signal_4456, signal_1622}), .b ({signal_5460, signal_5459, signal_5458, signal_1956}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({signal_5769, signal_5768, signal_5767, signal_2059}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2045 ( .a ({signal_4191, signal_4190, signal_4189, signal_1533}), .b ({signal_5475, signal_5474, signal_5473, signal_1961}), .clk ( clk ), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_5772, signal_5771, signal_5770, signal_2060}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2064 ( .a ({signal_5718, signal_5717, signal_5716, signal_2042}), .b ({signal_5829, signal_5828, signal_5827, signal_2079}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2068 ( .a ({signal_5733, signal_5732, signal_5731, signal_2047}), .b ({signal_5841, signal_5840, signal_5839, signal_2083}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2072 ( .a ({signal_5748, signal_5747, signal_5746, signal_2052}), .b ({signal_5853, signal_5852, signal_5851, signal_2087}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2073 ( .a ({signal_5766, signal_5765, signal_5764, signal_2058}), .b ({signal_5856, signal_5855, signal_5854, signal_2088}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2084 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_5544, signal_5543, signal_5542, signal_1984}), .clk ( clk ), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({signal_5889, signal_5888, signal_5887, signal_2099}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2090 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_5571, signal_5570, signal_5569, signal_1993}), .clk ( clk ), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({signal_5907, signal_5906, signal_5905, signal_2105}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2098 ( .a ({signal_5391, signal_5390, signal_5389, signal_1933}), .b ({signal_5589, signal_5588, signal_5587, signal_1999}), .clk ( clk ), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({signal_5931, signal_5930, signal_5929, signal_2113}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2100 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_5595, signal_5594, signal_5593, signal_2001}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({signal_5937, signal_5936, signal_5935, signal_2115}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2102 ( .a ({signal_5025, signal_5024, signal_5023, signal_1811}), .b ({signal_5604, signal_5603, signal_5602, signal_2004}), .clk ( clk ), .r ({Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_5943, signal_5942, signal_5941, signal_2117}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2103 ( .a ({signal_5532, signal_5531, signal_5530, signal_1980}), .b ({signal_5415, signal_5414, signal_5413, signal_1941}), .clk ( clk ), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086]}), .c ({signal_5946, signal_5945, signal_5944, signal_2118}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2105 ( .a ({signal_5541, signal_5540, signal_5539, signal_1983}), .b ({signal_5415, signal_5414, signal_5413, signal_1941}), .clk ( clk ), .r ({Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({signal_5952, signal_5951, signal_5950, signal_2120}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2106 ( .a ({signal_4365, signal_4364, signal_4363, signal_1591}), .b ({signal_5712, signal_5711, signal_5710, signal_2040}), .clk ( clk ), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098]}), .c ({signal_5955, signal_5954, signal_5953, signal_2121}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2107 ( .a ({signal_5487, signal_5486, signal_5485, signal_1965}), .b ({signal_5424, signal_5423, signal_5422, signal_1944}), .clk ( clk ), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({signal_5958, signal_5957, signal_5956, signal_2122}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2108 ( .a ({signal_5496, signal_5495, signal_5494, signal_1968}), .b ({signal_5727, signal_5726, signal_5725, signal_2045}), .clk ( clk ), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({signal_5961, signal_5960, signal_5959, signal_2123}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2109 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_5613, signal_5612, signal_5611, signal_2007}), .clk ( clk ), .r ({Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({signal_5964, signal_5963, signal_5962, signal_2124}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2111 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_5616, signal_5615, signal_5614, signal_2008}), .clk ( clk ), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122]}), .c ({signal_5970, signal_5969, signal_5968, signal_2126}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2112 ( .a ({signal_5502, signal_5501, signal_5500, signal_1970}), .b ({signal_5448, signal_5447, signal_5446, signal_1952}), .clk ( clk ), .r ({Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({signal_5973, signal_5972, signal_5971, signal_2127}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2113 ( .a ({signal_4455, signal_4454, signal_4453, signal_1621}), .b ({signal_5739, signal_5738, signal_5737, signal_2049}), .clk ( clk ), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134]}), .c ({signal_5976, signal_5975, signal_5974, signal_2128}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2114 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_5619, signal_5618, signal_5617, signal_2009}), .clk ( clk ), .r ({Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({signal_5979, signal_5978, signal_5977, signal_2129}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2115 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_5622, signal_5621, signal_5620, signal_2010}), .clk ( clk ), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146]}), .c ({signal_5982, signal_5981, signal_5980, signal_2130}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2117 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_5628, signal_5627, signal_5626, signal_2012}), .clk ( clk ), .r ({Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({signal_5988, signal_5987, signal_5986, signal_2132}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2120 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_5631, signal_5630, signal_5629, signal_2013}), .clk ( clk ), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158]}), .c ({signal_5997, signal_5996, signal_5995, signal_2135}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2129 ( .a ({signal_5889, signal_5888, signal_5887, signal_2099}), .b ({signal_6024, signal_6023, signal_6022, signal_2144}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2131 ( .a ({signal_5907, signal_5906, signal_5905, signal_2105}), .b ({signal_6030, signal_6029, signal_6028, signal_2146}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2132 ( .a ({signal_5937, signal_5936, signal_5935, signal_2115}), .b ({signal_6033, signal_6032, signal_6031, signal_2147}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2134 ( .a ({signal_5964, signal_5963, signal_5962, signal_2124}), .b ({signal_6039, signal_6038, signal_6037, signal_2149}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2136 ( .a ({signal_5970, signal_5969, signal_5968, signal_2126}), .b ({signal_6045, signal_6044, signal_6043, signal_2151}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2137 ( .a ({signal_5979, signal_5978, signal_5977, signal_2129}), .b ({signal_6048, signal_6047, signal_6046, signal_2152}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2138 ( .a ({signal_5982, signal_5981, signal_5980, signal_2130}), .b ({signal_6051, signal_6050, signal_6049, signal_2153}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2139 ( .a ({signal_5988, signal_5987, signal_5986, signal_2132}), .b ({signal_6054, signal_6053, signal_6052, signal_2154}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2141 ( .a ({signal_5997, signal_5996, signal_5995, signal_2135}), .b ({signal_6060, signal_6059, signal_6058, signal_2156}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2142 ( .a ({signal_3486, signal_3485, signal_3484, signal_1298}), .b ({signal_5775, signal_5774, signal_5773, signal_2061}), .clk ( clk ), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({signal_6063, signal_6062, signal_6061, signal_2157}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2143 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_5778, signal_5777, signal_5776, signal_2062}), .clk ( clk ), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({signal_6066, signal_6065, signal_6064, signal_2158}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2145 ( .a ({signal_4857, signal_4856, signal_4855, signal_1755}), .b ({signal_5862, signal_5861, signal_5860, signal_2090}), .clk ( clk ), .r ({Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({signal_6072, signal_6071, signal_6070, signal_2160}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2146 ( .a ({signal_5787, signal_5786, signal_5785, signal_2065}), .b ({signal_5553, signal_5552, signal_5551, signal_1987}), .clk ( clk ), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182]}), .c ({signal_6075, signal_6074, signal_6073, signal_2161}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2147 ( .a ({signal_4410, signal_4409, signal_4408, signal_1606}), .b ({signal_5790, signal_5789, signal_5788, signal_2066}), .clk ( clk ), .r ({Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({signal_6078, signal_6077, signal_6076, signal_2162}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2149 ( .a ({signal_4665, signal_4664, signal_4663, signal_1691}), .b ({signal_5871, signal_5870, signal_5869, signal_2093}), .clk ( clk ), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194]}), .c ({signal_6084, signal_6083, signal_6082, signal_2164}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2150 ( .a ({signal_4302, signal_4301, signal_4300, signal_1570}), .b ({signal_5874, signal_5873, signal_5872, signal_2094}), .clk ( clk ), .r ({Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({signal_6087, signal_6086, signal_6085, signal_2165}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2151 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_5808, signal_5807, signal_5806, signal_2072}), .clk ( clk ), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206]}), .c ({signal_6090, signal_6089, signal_6088, signal_2166}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2152 ( .a ({signal_2784, signal_2783, signal_2782, signal_1064}), .b ({signal_5877, signal_5876, signal_5875, signal_2095}), .clk ( clk ), .r ({Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({signal_6093, signal_6092, signal_6091, signal_2167}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2153 ( .a ({signal_4344, signal_4343, signal_4342, signal_1584}), .b ({signal_5886, signal_5885, signal_5884, signal_2098}), .clk ( clk ), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218]}), .c ({signal_6096, signal_6095, signal_6094, signal_2168}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2154 ( .a ({signal_3540, signal_3539, signal_3538, signal_1316}), .b ({signal_5817, signal_5816, signal_5815, signal_2075}), .clk ( clk ), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({signal_6099, signal_6098, signal_6097, signal_2169}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2155 ( .a ({signal_5784, signal_5783, signal_5782, signal_2064}), .b ({signal_5820, signal_5819, signal_5818, signal_2076}), .clk ( clk ), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({signal_6102, signal_6101, signal_6100, signal_2170}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2156 ( .a ({signal_4362, signal_4361, signal_4360, signal_1590}), .b ({signal_5823, signal_5822, signal_5821, signal_2077}), .clk ( clk ), .r ({Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({signal_6105, signal_6104, signal_6103, signal_2171}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2157 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_5826, signal_5825, signal_5824, signal_2078}), .clk ( clk ), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242]}), .c ({signal_6108, signal_6107, signal_6106, signal_2172}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2158 ( .a ({signal_4617, signal_4616, signal_4615, signal_1675}), .b ({signal_5892, signal_5891, signal_5890, signal_2100}), .clk ( clk ), .r ({Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({signal_6111, signal_6110, signal_6109, signal_2173}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2159 ( .a ({signal_4386, signal_4385, signal_4384, signal_1598}), .b ({signal_5898, signal_5897, signal_5896, signal_2102}), .clk ( clk ), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254]}), .c ({signal_6114, signal_6113, signal_6112, signal_2174}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2160 ( .a ({signal_5490, signal_5489, signal_5488, signal_1966}), .b ({signal_5901, signal_5900, signal_5899, signal_2103}), .clk ( clk ), .r ({Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({signal_6117, signal_6116, signal_6115, signal_2175}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2161 ( .a ({signal_4395, signal_4394, signal_4393, signal_1601}), .b ({signal_5904, signal_5903, signal_5902, signal_2104}), .clk ( clk ), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266]}), .c ({signal_6120, signal_6119, signal_6118, signal_2176}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2163 ( .a ({signal_4221, signal_4220, signal_4219, signal_1543}), .b ({signal_5832, signal_5831, signal_5830, signal_2080}), .clk ( clk ), .r ({Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({signal_6126, signal_6125, signal_6124, signal_2178}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2164 ( .a ({signal_3459, signal_3458, signal_3457, signal_1289}), .b ({signal_5913, signal_5912, signal_5911, signal_2107}), .clk ( clk ), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278]}), .c ({signal_6129, signal_6128, signal_6127, signal_2179}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2165 ( .a ({signal_5916, signal_5915, signal_5914, signal_2108}), .b ({signal_5451, signal_5450, signal_5449, signal_1953}), .clk ( clk ), .r ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284]}), .c ({signal_6132, signal_6131, signal_6130, signal_2180}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2166 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_5844, signal_5843, signal_5842, signal_2084}), .clk ( clk ), .r ({Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .c ({signal_6135, signal_6134, signal_6133, signal_2181}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2167 ( .a ({signal_5847, signal_5846, signal_5845, signal_2085}), .b ({signal_5625, signal_5624, signal_5623, signal_2011}), .clk ( clk ), .r ({Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296]}), .c ({signal_6138, signal_6137, signal_6136, signal_2182}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2168 ( .a ({signal_5121, signal_5120, signal_5119, signal_1843}), .b ({signal_5928, signal_5927, signal_5926, signal_2112}), .clk ( clk ), .r ({Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302]}), .c ({signal_6141, signal_6140, signal_6139, signal_2183}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2169 ( .a ({signal_4467, signal_4466, signal_4465, signal_1625}), .b ({signal_5850, signal_5849, signal_5848, signal_2086}), .clk ( clk ), .r ({Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308]}), .c ({signal_6144, signal_6143, signal_6142, signal_2184}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2171 ( .a ({signal_3669, signal_3668, signal_3667, signal_1359}), .b ({signal_5934, signal_5933, signal_5932, signal_2114}), .clk ( clk ), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314]}), .c ({signal_6150, signal_6149, signal_6148, signal_2186}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2184 ( .a ({signal_6066, signal_6065, signal_6064, signal_2158}), .b ({signal_6189, signal_6188, signal_6187, signal_2199}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2187 ( .a ({signal_6090, signal_6089, signal_6088, signal_2166}), .b ({signal_6198, signal_6197, signal_6196, signal_2202}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2188 ( .a ({signal_6108, signal_6107, signal_6106, signal_2172}), .b ({signal_6201, signal_6200, signal_6199, signal_2203}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2189 ( .a ({signal_6114, signal_6113, signal_6112, signal_2174}), .b ({signal_6204, signal_6203, signal_6202, signal_2204}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2191 ( .a ({signal_6129, signal_6128, signal_6127, signal_2179}), .b ({signal_6210, signal_6209, signal_6208, signal_2206}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2192 ( .a ({signal_6132, signal_6131, signal_6130, signal_2180}), .b ({signal_6213, signal_6212, signal_6211, signal_2207}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2193 ( .a ({signal_6135, signal_6134, signal_6133, signal_2181}), .b ({signal_6216, signal_6215, signal_6214, signal_2208}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2194 ( .a ({signal_6150, signal_6149, signal_6148, signal_2186}), .b ({signal_6219, signal_6218, signal_6217, signal_2209}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2201 ( .a ({signal_3513, signal_3512, signal_3511, signal_1307}), .b ({signal_6009, signal_6008, signal_6007, signal_2139}), .clk ( clk ), .r ({Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({signal_6240, signal_6239, signal_6238, signal_2216}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2202 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_6012, signal_6011, signal_6010, signal_2140}), .clk ( clk ), .r ({Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326]}), .c ({signal_6243, signal_6242, signal_6241, signal_2217}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2203 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_6015, signal_6014, signal_6013, signal_2141}), .clk ( clk ), .r ({Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332]}), .c ({signal_6246, signal_6245, signal_6244, signal_2218}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2204 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_6018, signal_6017, signal_6016, signal_2142}), .clk ( clk ), .r ({Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338]}), .c ({signal_6249, signal_6248, signal_6247, signal_2219}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2205 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_6021, signal_6020, signal_6019, signal_2143}), .clk ( clk ), .r ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344]}), .c ({signal_6252, signal_6251, signal_6250, signal_2220}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2206 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_6027, signal_6026, signal_6025, signal_2145}), .clk ( clk ), .r ({Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .c ({signal_6255, signal_6254, signal_6253, signal_2221}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2213 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_6036, signal_6035, signal_6034, signal_2148}), .clk ( clk ), .r ({Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356]}), .c ({signal_6276, signal_6275, signal_6274, signal_2228}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2221 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_6042, signal_6041, signal_6040, signal_2150}), .clk ( clk ), .r ({Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362]}), .c ({signal_6300, signal_6299, signal_6298, signal_2236}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2233 ( .a ({signal_6240, signal_6239, signal_6238, signal_2216}), .b ({signal_6336, signal_6335, signal_6334, signal_2248}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2234 ( .a ({signal_6243, signal_6242, signal_6241, signal_2217}), .b ({signal_6339, signal_6338, signal_6337, signal_2249}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2235 ( .a ({signal_6246, signal_6245, signal_6244, signal_2218}), .b ({signal_6342, signal_6341, signal_6340, signal_2250}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2236 ( .a ({signal_6249, signal_6248, signal_6247, signal_2219}), .b ({signal_6345, signal_6344, signal_6343, signal_2251}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2237 ( .a ({signal_6252, signal_6251, signal_6250, signal_2220}), .b ({signal_6348, signal_6347, signal_6346, signal_2252}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2238 ( .a ({signal_6255, signal_6254, signal_6253, signal_2221}), .b ({signal_6351, signal_6350, signal_6349, signal_2253}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2240 ( .a ({signal_6276, signal_6275, signal_6274, signal_2228}), .b ({signal_6357, signal_6356, signal_6355, signal_2255}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2242 ( .a ({signal_6300, signal_6299, signal_6298, signal_2236}), .b ({signal_6363, signal_6362, signal_6361, signal_2257}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2248 ( .a ({signal_5814, signal_5813, signal_5812, signal_2074}), .b ({signal_6192, signal_6191, signal_6190, signal_2200}), .clk ( clk ), .r ({Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368]}), .c ({signal_6381, signal_6380, signal_6379, signal_2263}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2116 ( .a ({signal_3537, signal_3536, signal_3535, signal_1315}), .b ({signal_5751, signal_5750, signal_5749, signal_2053}), .clk ( clk ), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374]}), .c ({signal_5985, signal_5984, signal_5983, signal_2131}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2118 ( .a ({signal_4866, signal_4865, signal_4864, signal_1758}), .b ({signal_5754, signal_5753, signal_5752, signal_2054}), .clk ( clk ), .r ({Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({signal_5991, signal_5990, signal_5989, signal_2133}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2119 ( .a ({signal_4527, signal_4526, signal_4525, signal_1645}), .b ({signal_5757, signal_5756, signal_5755, signal_2055}), .clk ( clk ), .r ({Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386]}), .c ({signal_5994, signal_5993, signal_5992, signal_2134}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2121 ( .a ({signal_4440, signal_4439, signal_4438, signal_1616}), .b ({signal_5763, signal_5762, signal_5761, signal_2057}), .clk ( clk ), .r ({Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392]}), .c ({signal_6000, signal_5999, signal_5998, signal_2136}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2122 ( .a ({signal_4878, signal_4877, signal_4876, signal_1762}), .b ({signal_5769, signal_5768, signal_5767, signal_2059}), .clk ( clk ), .r ({Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398]}), .c ({signal_6003, signal_6002, signal_6001, signal_2137}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2123 ( .a ({signal_4194, signal_4193, signal_4192, signal_1534}), .b ({signal_5772, signal_5771, signal_5770, signal_2060}), .clk ( clk ), .r ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404]}), .c ({signal_6006, signal_6005, signal_6004, signal_2138}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2140 ( .a ({signal_5994, signal_5993, signal_5992, signal_2134}), .b ({signal_6057, signal_6056, signal_6055, signal_2155}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2162 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_5829, signal_5828, signal_5827, signal_2079}), .clk ( clk ), .r ({Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .c ({signal_6123, signal_6122, signal_6121, signal_2177}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2170 ( .a ({signal_5127, signal_5126, signal_5125, signal_1845}), .b ({signal_5931, signal_5930, signal_5929, signal_2113}), .clk ( clk ), .r ({Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416]}), .c ({signal_6147, signal_6146, signal_6145, signal_2185}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2172 ( .a ({signal_5805, signal_5804, signal_5803, signal_2071}), .b ({signal_5943, signal_5942, signal_5941, signal_2117}), .clk ( clk ), .r ({Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422]}), .c ({signal_6153, signal_6152, signal_6151, signal_2187}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2173 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_5853, signal_5852, signal_5851, signal_2087}), .clk ( clk ), .r ({Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428]}), .c ({signal_6156, signal_6155, signal_6154, signal_2188}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2174 ( .a ({signal_5142, signal_5141, signal_5140, signal_1850}), .b ({signal_5955, signal_5954, signal_5953, signal_2121}), .clk ( clk ), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434]}), .c ({signal_6159, signal_6158, signal_6157, signal_2189}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2175 ( .a ({signal_4485, signal_4484, signal_4483, signal_1631}), .b ({signal_5958, signal_5957, signal_5956, signal_2122}), .clk ( clk ), .r ({Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({signal_6162, signal_6161, signal_6160, signal_2190}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2176 ( .a ({signal_4641, signal_4640, signal_4639, signal_1683}), .b ({signal_5961, signal_5960, signal_5959, signal_2123}), .clk ( clk ), .r ({Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446]}), .c ({signal_6165, signal_6164, signal_6163, signal_2191}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2177 ( .a ({signal_5841, signal_5840, signal_5839, signal_2083}), .b ({signal_5760, signal_5759, signal_5758, signal_2056}), .clk ( clk ), .r ({Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452]}), .c ({signal_6168, signal_6167, signal_6166, signal_2192}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2178 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_5856, signal_5855, signal_5854, signal_2088}), .clk ( clk ), .r ({Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458]}), .c ({signal_6171, signal_6170, signal_6169, signal_2193}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2179 ( .a ({signal_5022, signal_5021, signal_5020, signal_1810}), .b ({signal_5976, signal_5975, signal_5974, signal_2128}), .clk ( clk ), .r ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464]}), .c ({signal_6174, signal_6173, signal_6172, signal_2194}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2190 ( .a ({signal_6123, signal_6122, signal_6121, signal_2177}), .b ({signal_6207, signal_6206, signal_6205, signal_2205}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2195 ( .a ({signal_6156, signal_6155, signal_6154, signal_2188}), .b ({signal_6222, signal_6221, signal_6220, signal_2210}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2196 ( .a ({signal_6162, signal_6161, signal_6160, signal_2190}), .b ({signal_6225, signal_6224, signal_6223, signal_2211}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2197 ( .a ({signal_6165, signal_6164, signal_6163, signal_2191}), .b ({signal_6228, signal_6227, signal_6226, signal_2212}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2198 ( .a ({signal_6171, signal_6170, signal_6169, signal_2193}), .b ({signal_6231, signal_6230, signal_6229, signal_2213}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2200 ( .a ({signal_3489, signal_3488, signal_3487, signal_1299}), .b ({signal_6063, signal_6062, signal_6061, signal_2157}), .clk ( clk ), .r ({Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .c ({signal_6237, signal_6236, signal_6235, signal_2215}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2207 ( .a ({signal_5835, signal_5834, signal_5833, signal_2081}), .b ({signal_6030, signal_6029, signal_6028, signal_2146}), .clk ( clk ), .r ({Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476]}), .c ({signal_6258, signal_6257, signal_6256, signal_2222}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2208 ( .a ({signal_4263, signal_4262, signal_4261, signal_1557}), .b ({signal_6084, signal_6083, signal_6082, signal_2164}), .clk ( clk ), .r ({Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482]}), .c ({signal_6261, signal_6260, signal_6259, signal_2223}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2209 ( .a ({signal_5799, signal_5798, signal_5797, signal_2069}), .b ({signal_6033, signal_6032, signal_6031, signal_2147}), .clk ( clk ), .r ({Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488]}), .c ({signal_6264, signal_6263, signal_6262, signal_2224}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2210 ( .a ({signal_3309, signal_3308, signal_3307, signal_1239}), .b ({signal_6087, signal_6086, signal_6085, signal_2165}), .clk ( clk ), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494]}), .c ({signal_6267, signal_6266, signal_6265, signal_2225}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2211 ( .a ({signal_5034, signal_5033, signal_5032, signal_1814}), .b ({signal_6093, signal_6092, signal_6091, signal_2167}), .clk ( clk ), .r ({Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({signal_6270, signal_6269, signal_6268, signal_2226}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2212 ( .a ({signal_5946, signal_5945, signal_5944, signal_2118}), .b ({signal_6096, signal_6095, signal_6094, signal_2168}), .clk ( clk ), .r ({Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506]}), .c ({signal_6273, signal_6272, signal_6271, signal_2227}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2214 ( .a ({signal_5052, signal_5051, signal_5050, signal_1820}), .b ({signal_6099, signal_6098, signal_6097, signal_2169}), .clk ( clk ), .r ({Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512]}), .c ({signal_6279, signal_6278, signal_6277, signal_2229}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2215 ( .a ({signal_5952, signal_5951, signal_5950, signal_2120}), .b ({signal_6102, signal_6101, signal_6100, signal_2170}), .clk ( clk ), .r ({Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518]}), .c ({signal_6282, signal_6281, signal_6280, signal_2230}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2216 ( .a ({signal_4110, signal_4109, signal_4108, signal_1506}), .b ({signal_6105, signal_6104, signal_6103, signal_2171}), .clk ( clk ), .r ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524]}), .c ({signal_6285, signal_6284, signal_6283, signal_2231}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2217 ( .a ({signal_4371, signal_4370, signal_4369, signal_1593}), .b ({signal_6111, signal_6110, signal_6109, signal_2173}), .clk ( clk ), .r ({Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .c ({signal_6288, signal_6287, signal_6286, signal_2232}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2218 ( .a ({signal_5610, signal_5609, signal_5608, signal_2006}), .b ({signal_6117, signal_6116, signal_6115, signal_2175}), .clk ( clk ), .r ({Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536]}), .c ({signal_6291, signal_6290, signal_6289, signal_2233}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2219 ( .a ({signal_2772, signal_2771, signal_2770, signal_1060}), .b ({signal_6120, signal_6119, signal_6118, signal_2176}), .clk ( clk ), .r ({Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542]}), .c ({signal_6294, signal_6293, signal_6292, signal_2234}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2220 ( .a ({signal_3606, signal_3605, signal_3604, signal_1338}), .b ({signal_6126, signal_6125, signal_6124, signal_2178}), .clk ( clk ), .r ({Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548]}), .c ({signal_6297, signal_6296, signal_6295, signal_2235}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2222 ( .a ({signal_6045, signal_6044, signal_6043, signal_2151}), .b ({signal_5973, signal_5972, signal_5971, signal_2127}), .clk ( clk ), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554]}), .c ({signal_6303, signal_6302, signal_6301, signal_2237}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2223 ( .a ({signal_6051, signal_6050, signal_6049, signal_2153}), .b ({signal_6138, signal_6137, signal_6136, signal_2182}), .clk ( clk ), .r ({Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({signal_6306, signal_6305, signal_6304, signal_2238}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2224 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_6144, signal_6143, signal_6142, signal_2184}), .clk ( clk ), .r ({Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566]}), .c ({signal_6309, signal_6308, signal_6307, signal_2239}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2239 ( .a ({signal_6261, signal_6260, signal_6259, signal_2223}), .b ({signal_6354, signal_6353, signal_6352, signal_2254}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2241 ( .a ({signal_6288, signal_6287, signal_6286, signal_2232}), .b ({signal_6360, signal_6359, signal_6358, signal_2256}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2243 ( .a ({signal_6309, signal_6308, signal_6307, signal_2239}), .b ({signal_6366, signal_6365, signal_6364, signal_2258}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2249 ( .a ({signal_6078, signal_6077, signal_6076, signal_2162}), .b ({signal_6195, signal_6194, signal_6193, signal_2201}), .clk ( clk ), .r ({Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572]}), .c ({signal_6384, signal_6383, signal_6382, signal_2264}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2250 ( .a ({signal_6024, signal_6023, signal_6022, signal_2144}), .b ({signal_6201, signal_6200, signal_6199, signal_2203}), .clk ( clk ), .r ({Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578]}), .c ({signal_6387, signal_6386, signal_6385, signal_2265}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2251 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_6204, signal_6203, signal_6202, signal_2204}), .clk ( clk ), .r ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584]}), .c ({signal_6390, signal_6389, signal_6388, signal_2266}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2252 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_6210, signal_6209, signal_6208, signal_2206}), .clk ( clk ), .r ({Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .c ({signal_6393, signal_6392, signal_6391, signal_2267}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2253 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_6213, signal_6212, signal_6211, signal_2207}), .clk ( clk ), .r ({Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596]}), .c ({signal_6396, signal_6395, signal_6394, signal_2268}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2254 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_6219, signal_6218, signal_6217, signal_2209}), .clk ( clk ), .r ({Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602]}), .c ({signal_6399, signal_6398, signal_6397, signal_2269}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2271 ( .a ({signal_6390, signal_6389, signal_6388, signal_2266}), .b ({signal_6450, signal_6449, signal_6448, signal_2286}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2272 ( .a ({signal_6393, signal_6392, signal_6391, signal_2267}), .b ({signal_6453, signal_6452, signal_6451, signal_2287}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2273 ( .a ({signal_6396, signal_6395, signal_6394, signal_2268}), .b ({signal_6456, signal_6455, signal_6454, signal_2288}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2274 ( .a ({signal_6399, signal_6398, signal_6397, signal_2269}), .b ({signal_6459, signal_6458, signal_6457, signal_2289}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2282 ( .a ({signal_6342, signal_6341, signal_6340, signal_2250}), .b ({signal_4503, signal_4502, signal_4501, signal_1637}), .clk ( clk ), .r ({Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608]}), .c ({signal_6483, signal_6482, signal_6481, signal_2297}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2283 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_6336, signal_6335, signal_6334, signal_2248}), .clk ( clk ), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614]}), .c ({signal_6486, signal_6485, signal_6484, signal_2298}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2285 ( .a ({signal_4146, signal_4145, signal_4144, signal_1518}), .b ({signal_6381, signal_6380, signal_6379, signal_2263}), .clk ( clk ), .r ({Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({signal_6492, signal_6491, signal_6490, signal_2300}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2286 ( .a ({signal_5046, signal_5045, signal_5044, signal_1818}), .b ({signal_6345, signal_6344, signal_6343, signal_2251}), .clk ( clk ), .r ({Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626]}), .c ({signal_6495, signal_6494, signal_6493, signal_2301}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2297 ( .a ({signal_6486, signal_6485, signal_6484, signal_2298}), .b ({signal_6528, signal_6527, signal_6526, signal_2312}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2180 ( .a ({signal_3354, signal_3353, signal_3352, signal_1254}), .b ({signal_5985, signal_5984, signal_5983, signal_2131}), .clk ( clk ), .r ({Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632]}), .c ({signal_6177, signal_6176, signal_6175, signal_2195}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2181 ( .a ({signal_5556, signal_5555, signal_5554, signal_1988}), .b ({signal_5991, signal_5990, signal_5989, signal_2133}), .clk ( clk ), .r ({Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638]}), .c ({signal_6180, signal_6179, signal_6178, signal_2196}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2182 ( .a ({signal_4449, signal_4448, signal_4447, signal_1619}), .b ({signal_6000, signal_5999, signal_5998, signal_2136}), .clk ( clk ), .r ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644]}), .c ({signal_6183, signal_6182, signal_6181, signal_2197}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2183 ( .a ({signal_3642, signal_3641, signal_3640, signal_1350}), .b ({signal_6003, signal_6002, signal_6001, signal_2137}), .clk ( clk ), .r ({Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .c ({signal_6186, signal_6185, signal_6184, signal_2198}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2199 ( .a ({signal_6177, signal_6176, signal_6175, signal_2195}), .b ({signal_6234, signal_6233, signal_6232, signal_2214}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2225 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_6147, signal_6146, signal_6145, signal_2185}), .clk ( clk ), .r ({Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656]}), .c ({signal_6312, signal_6311, signal_6310, signal_2240}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2226 ( .a ({signal_5940, signal_5939, signal_5938, signal_2116}), .b ({signal_6153, signal_6152, signal_6151, signal_2187}), .clk ( clk ), .r ({Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662]}), .c ({signal_6315, signal_6314, signal_6313, signal_2241}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2227 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_6057, signal_6056, signal_6055, signal_2155}), .clk ( clk ), .r ({Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668]}), .c ({signal_6318, signal_6317, signal_6316, signal_2242}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2228 ( .a ({signal_6168, signal_6167, signal_6166, signal_2192}), .b ({signal_6060, signal_6059, signal_6058, signal_2156}), .clk ( clk ), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674]}), .c ({signal_6321, signal_6320, signal_6319, signal_2243}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2229 ( .a ({signal_5919, signal_5918, signal_5917, signal_2109}), .b ({signal_6174, signal_6173, signal_6172, signal_2194}), .clk ( clk ), .r ({Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({signal_6324, signal_6323, signal_6322, signal_2244}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2244 ( .a ({signal_6312, signal_6311, signal_6310, signal_2240}), .b ({signal_6369, signal_6368, signal_6367, signal_2259}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2245 ( .a ({signal_6318, signal_6317, signal_6316, signal_2242}), .b ({signal_6372, signal_6371, signal_6370, signal_2260}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2246 ( .a ({signal_6324, signal_6323, signal_6322, signal_2244}), .b ({signal_6375, signal_6374, signal_6373, signal_2261}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2247 ( .a ({signal_3333, signal_3332, signal_3331, signal_1247}), .b ({signal_6237, signal_6236, signal_6235, signal_2215}), .clk ( clk ), .r ({Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686]}), .c ({signal_6378, signal_6377, signal_6376, signal_2262}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2255 ( .a ({signal_5640, signal_5639, signal_5638, signal_2016}), .b ({signal_6264, signal_6263, signal_6262, signal_2224}), .clk ( clk ), .r ({Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692]}), .c ({signal_6402, signal_6401, signal_6400, signal_2270}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2256 ( .a ({signal_5022, signal_5021, signal_5020, signal_1810}), .b ({signal_6267, signal_6266, signal_6265, signal_2225}), .clk ( clk ), .r ({Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698]}), .c ({signal_6405, signal_6404, signal_6403, signal_2271}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2257 ( .a ({signal_4317, signal_4316, signal_4315, signal_1575}), .b ({signal_6270, signal_6269, signal_6268, signal_2226}), .clk ( clk ), .r ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704]}), .c ({signal_6408, signal_6407, signal_6406, signal_2272}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2258 ( .a ({signal_5529, signal_5528, signal_5527, signal_1979}), .b ({signal_6273, signal_6272, signal_6271, signal_2227}), .clk ( clk ), .r ({Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .c ({signal_6411, signal_6410, signal_6409, signal_2273}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2259 ( .a ({signal_4353, signal_4352, signal_4351, signal_1587}), .b ({signal_6279, signal_6278, signal_6277, signal_2229}), .clk ( clk ), .r ({Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716]}), .c ({signal_6414, signal_6413, signal_6412, signal_2274}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2260 ( .a ({signal_5175, signal_5174, signal_5173, signal_1861}), .b ({signal_6282, signal_6281, signal_6280, signal_2230}), .clk ( clk ), .r ({Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722]}), .c ({signal_6417, signal_6416, signal_6415, signal_2275}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2261 ( .a ({signal_3366, signal_3365, signal_3364, signal_1258}), .b ({signal_6285, signal_6284, signal_6283, signal_2231}), .clk ( clk ), .r ({Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728]}), .c ({signal_6420, signal_6419, signal_6418, signal_2276}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2262 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_6225, signal_6224, signal_6223, signal_2211}), .clk ( clk ), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734]}), .c ({signal_6423, signal_6422, signal_6421, signal_2277}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2263 ( .a ({signal_2790, signal_2789, signal_2788, signal_1066}), .b ({signal_6294, signal_6293, signal_6292, signal_2234}), .clk ( clk ), .r ({Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({signal_6426, signal_6425, signal_6424, signal_2278}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2264 ( .a ({signal_6207, signal_6206, signal_6205, signal_2205}), .b ({signal_6297, signal_6296, signal_6295, signal_2235}), .clk ( clk ), .r ({Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746]}), .c ({signal_6429, signal_6428, signal_6427, signal_2279}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2265 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_6228, signal_6227, signal_6226, signal_2212}), .clk ( clk ), .r ({Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752]}), .c ({signal_6432, signal_6431, signal_6430, signal_2280}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2266 ( .a ({signal_4434, signal_4433, signal_4432, signal_1614}), .b ({signal_6303, signal_6302, signal_6301, signal_2237}), .clk ( clk ), .r ({Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758]}), .c ({signal_6435, signal_6434, signal_6433, signal_2281}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2275 ( .a ({signal_6405, signal_6404, signal_6403, signal_2271}), .b ({signal_6462, signal_6461, signal_6460, signal_2290}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2276 ( .a ({signal_6408, signal_6407, signal_6406, signal_2272}), .b ({signal_6465, signal_6464, signal_6463, signal_2291}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2277 ( .a ({signal_6414, signal_6413, signal_6412, signal_2274}), .b ({signal_6468, signal_6467, signal_6466, signal_2292}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2278 ( .a ({signal_6420, signal_6419, signal_6418, signal_2276}), .b ({signal_6471, signal_6470, signal_6469, signal_2293}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2279 ( .a ({signal_6423, signal_6422, signal_6421, signal_2277}), .b ({signal_6474, signal_6473, signal_6472, signal_2294}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2280 ( .a ({signal_6432, signal_6431, signal_6430, signal_2280}), .b ({signal_6477, signal_6476, signal_6475, signal_2295}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2287 ( .a ({signal_6384, signal_6383, signal_6382, signal_2264}), .b ({signal_6258, signal_6257, signal_6256, signal_2222}), .clk ( clk ), .r ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764]}), .c ({signal_6498, signal_6497, signal_6496, signal_2302}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2288 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_6354, signal_6353, signal_6352, signal_2254}), .clk ( clk ), .r ({Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .c ({signal_6501, signal_6500, signal_6499, signal_2303}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2290 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_6360, signal_6359, signal_6358, signal_2256}), .clk ( clk ), .r ({Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776]}), .c ({signal_6507, signal_6506, signal_6505, signal_2305}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2299 ( .a ({signal_6501, signal_6500, signal_6499, signal_2303}), .b ({signal_6534, signal_6533, signal_6532, signal_2314}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2301 ( .a ({signal_6507, signal_6506, signal_6505, signal_2305}), .b ({signal_6540, signal_6539, signal_6538, signal_2316}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2304 ( .a ({signal_4239, signal_4238, signal_4237, signal_1549}), .b ({signal_6483, signal_6482, signal_6481, signal_2297}), .clk ( clk ), .r ({Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782]}), .c ({signal_6549, signal_6548, signal_6547, signal_2319}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2305 ( .a ({signal_4326, signal_4325, signal_4324, signal_1578}), .b ({signal_6492, signal_6491, signal_6490, signal_2300}), .clk ( clk ), .r ({Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788]}), .c ({signal_6552, signal_6551, signal_6550, signal_2320}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2306 ( .a ({signal_4335, signal_4334, signal_4333, signal_1581}), .b ({signal_6495, signal_6494, signal_6493, signal_2301}), .clk ( clk ), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794]}), .c ({signal_6555, signal_6554, signal_6553, signal_2321}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2307 ( .a ({signal_6450, signal_6449, signal_6448, signal_2286}), .b ({signal_6291, signal_6290, signal_6289, signal_2233}), .clk ( clk ), .r ({Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({signal_6558, signal_6557, signal_6556, signal_2322}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2230 ( .a ({signal_5427, signal_5426, signal_5425, signal_1945}), .b ({signal_6180, signal_6179, signal_6178, signal_2196}), .clk ( clk ), .r ({Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806]}), .c ({signal_6327, signal_6326, signal_6325, signal_2245}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2231 ( .a ({signal_5682, signal_5681, signal_5680, signal_2030}), .b ({signal_6183, signal_6182, signal_6181, signal_2197}), .clk ( clk ), .r ({Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812]}), .c ({signal_6330, signal_6329, signal_6328, signal_2246}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2232 ( .a ({signal_5925, signal_5924, signal_5923, signal_2111}), .b ({signal_6186, signal_6185, signal_6184, signal_2198}), .clk ( clk ), .r ({Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818]}), .c ({signal_6333, signal_6332, signal_6331, signal_2247}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2267 ( .a ({signal_5520, signal_5519, signal_5518, signal_1976}), .b ({signal_6315, signal_6314, signal_6313, signal_2241}), .clk ( clk ), .r ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824]}), .c ({signal_6438, signal_6437, signal_6436, signal_2282}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2268 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_6234, signal_6233, signal_6232, signal_2214}), .clk ( clk ), .r ({Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .c ({signal_6441, signal_6440, signal_6439, signal_2283}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2281 ( .a ({signal_6441, signal_6440, signal_6439, signal_2283}), .b ({signal_6480, signal_6479, signal_6478, signal_2296}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2284 ( .a ({signal_4107, signal_4106, signal_4105, signal_1505}), .b ({signal_6378, signal_6377, signal_6376, signal_2262}), .clk ( clk ), .r ({Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836]}), .c ({signal_6489, signal_6488, signal_6487, signal_2299}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2289 ( .a ({signal_6366, signal_6365, signal_6364, signal_2258}), .b ({signal_6369, signal_6368, signal_6367, signal_2259}), .clk ( clk ), .r ({Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842]}), .c ({signal_6504, signal_6503, signal_6502, signal_2304}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2291 ( .a ({signal_5802, signal_5801, signal_5800, signal_2070}), .b ({signal_6402, signal_6401, signal_6400, signal_2270}), .clk ( clk ), .r ({Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848]}), .c ({signal_6510, signal_6509, signal_6508, signal_2306}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2292 ( .a ({signal_5538, signal_5537, signal_5536, signal_1982}), .b ({signal_6411, signal_6410, signal_6409, signal_2273}), .clk ( clk ), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854]}), .c ({signal_6513, signal_6512, signal_6511, signal_2307}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2293 ( .a ({signal_4359, signal_4358, signal_4357, signal_1589}), .b ({signal_6417, signal_6416, signal_6415, signal_2275}), .clk ( clk ), .r ({Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({signal_6516, signal_6515, signal_6514, signal_2308}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2294 ( .a ({signal_5493, signal_5492, signal_5491, signal_1967}), .b ({signal_6426, signal_6425, signal_6424, signal_2278}), .clk ( clk ), .r ({Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866]}), .c ({signal_6519, signal_6518, signal_6517, signal_2309}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2295 ( .a ({signal_5262, signal_5261, signal_5260, signal_1890}), .b ({signal_6375, signal_6374, signal_6373, signal_2261}), .clk ( clk ), .r ({Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872]}), .c ({signal_6522, signal_6521, signal_6520, signal_2310}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2298 ( .a ({signal_6489, signal_6488, signal_6487, signal_2299}), .b ({signal_6531, signal_6530, signal_6529, signal_2313}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2300 ( .a ({signal_6504, signal_6503, signal_6502, signal_2304}), .b ({signal_6537, signal_6536, signal_6535, signal_2315}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2302 ( .a ({signal_6519, signal_6518, signal_6517, signal_2309}), .b ({signal_6543, signal_6542, signal_6541, signal_2317}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2303 ( .a ({signal_6522, signal_6521, signal_6520, signal_2310}), .b ({signal_6546, signal_6545, signal_6544, signal_2318}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2308 ( .a ({signal_5598, signal_5597, signal_5596, signal_2002}), .b ({signal_6462, signal_6461, signal_6460, signal_2290}), .clk ( clk ), .r ({Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878]}), .c ({signal_6561, signal_6560, signal_6559, signal_2323}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2309 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_6465, signal_6464, signal_6463, signal_2291}), .clk ( clk ), .r ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884]}), .c ({signal_6564, signal_6563, signal_6562, signal_2324}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2310 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_6468, signal_6467, signal_6466, signal_2292}), .clk ( clk ), .r ({Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .c ({signal_6567, signal_6566, signal_6565, signal_2325}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2311 ( .a ({signal_2439, signal_2438, signal_2437, signal_949}), .b ({signal_6471, signal_6470, signal_6469, signal_2293}), .clk ( clk ), .r ({Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896]}), .c ({signal_6570, signal_6569, signal_6568, signal_2326}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2312 ( .a ({signal_6351, signal_6350, signal_6349, signal_2253}), .b ({signal_6474, signal_6473, signal_6472, signal_2294}), .clk ( clk ), .r ({Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902]}), .c ({signal_6573, signal_6572, signal_6571, signal_2327}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2313 ( .a ({signal_6498, signal_6497, signal_6496, signal_2302}), .b ({signal_6429, signal_6428, signal_6427, signal_2279}), .clk ( clk ), .r ({Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908]}), .c ({signal_6576, signal_6575, signal_6574, signal_2328}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2314 ( .a ({signal_5910, signal_5909, signal_5908, signal_2106}), .b ({signal_6477, signal_6476, signal_6475, signal_2295}), .clk ( clk ), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914]}), .c ({signal_6579, signal_6578, signal_6577, signal_2329}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2315 ( .a ({signal_6453, signal_6452, signal_6451, signal_2287}), .b ({signal_6321, signal_6320, signal_6319, signal_2243}), .clk ( clk ), .r ({Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({signal_6582, signal_6581, signal_6580, signal_2330}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2320 ( .a ({signal_6561, signal_6560, signal_6559, signal_2323}), .b ({signal_6597, signal_6596, signal_6595, signal_2335}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2321 ( .a ({signal_6564, signal_6563, signal_6562, signal_2324}), .b ({signal_6600, signal_6599, signal_6598, signal_2336}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2322 ( .a ({signal_6567, signal_6566, signal_6565, signal_2325}), .b ({signal_6603, signal_6602, signal_6601, signal_2337}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2323 ( .a ({signal_6570, signal_6569, signal_6568, signal_2326}), .b ({signal_6606, signal_6605, signal_6604, signal_2338}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2324 ( .a ({signal_5796, signal_5795, signal_5794, signal_2068}), .b ({signal_6549, signal_6548, signal_6547, signal_2319}), .clk ( clk ), .r ({Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926]}), .c ({signal_6609, signal_6608, signal_6607, signal_2339}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2326 ( .a ({signal_6216, signal_6215, signal_6214, signal_2208}), .b ({signal_6534, signal_6533, signal_6532, signal_2314}), .clk ( clk ), .r ({Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932]}), .c ({signal_6615, signal_6614, signal_6613, signal_2341}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2328 ( .a ({signal_5811, signal_5810, signal_5809, signal_2073}), .b ({signal_6552, signal_6551, signal_6550, signal_2320}), .clk ( clk ), .r ({Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938]}), .c ({signal_6621, signal_6620, signal_6619, signal_2343}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2329 ( .a ({signal_6528, signal_6527, signal_6526, signal_2312}), .b ({signal_6555, signal_6554, signal_6553, signal_2321}), .clk ( clk ), .r ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944]}), .c ({signal_6624, signal_6623, signal_6622, signal_2344}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2330 ( .a ({signal_6339, signal_6338, signal_6337, signal_2249}), .b ({signal_6540, signal_6539, signal_6538, signal_2316}), .clk ( clk ), .r ({Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .c ({signal_6627, signal_6626, signal_6625, signal_2345}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2269 ( .a ({signal_6075, signal_6074, signal_6073, signal_2161}), .b ({signal_6327, signal_6326, signal_6325, signal_2245}), .clk ( clk ), .r ({Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956]}), .c ({signal_6444, signal_6443, signal_6442, signal_2284}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2270 ( .a ({signal_5922, signal_5921, signal_5920, signal_2110}), .b ({signal_6333, signal_6332, signal_6331, signal_2247}), .clk ( clk ), .r ({Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962]}), .c ({signal_6447, signal_6446, signal_6445, signal_2285}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2296 ( .a ({signal_6189, signal_6188, signal_6187, signal_2199}), .b ({signal_6438, signal_6437, signal_6436, signal_2282}), .clk ( clk ), .r ({Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968]}), .c ({signal_6525, signal_6524, signal_6523, signal_2311}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2316 ( .a ({signal_5526, signal_5525, signal_5524, signal_1978}), .b ({signal_6513, signal_6512, signal_6511, signal_2307}), .clk ( clk ), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974]}), .c ({signal_6585, signal_6584, signal_6583, signal_2331}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2317 ( .a ({signal_6357, signal_6356, signal_6355, signal_2255}), .b ({signal_6480, signal_6479, signal_6478, signal_2296}), .clk ( clk ), .r ({Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({signal_6588, signal_6587, signal_6586, signal_2332}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2318 ( .a ({signal_6456, signal_6455, signal_6454, signal_2288}), .b ({signal_6330, signal_6329, signal_6328, signal_2246}), .clk ( clk ), .r ({Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986]}), .c ({signal_6591, signal_6590, signal_6589, signal_2333}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2325 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_6531, signal_6530, signal_6529, signal_2313}), .clk ( clk ), .r ({Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992]}), .c ({signal_6612, signal_6611, signal_6610, signal_2340}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2327 ( .a ({signal_6141, signal_6140, signal_6139, signal_2183}), .b ({signal_6537, signal_6536, signal_6535, signal_2315}), .clk ( clk ), .r ({Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998]}), .c ({signal_6618, signal_6617, signal_6616, signal_2342}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2331 ( .a ({signal_5550, signal_5549, signal_5548, signal_1986}), .b ({signal_6573, signal_6572, signal_6571, signal_2327}), .clk ( clk ), .r ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004]}), .c ({signal_6630, signal_6629, signal_6628, signal_2346}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2332 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_6543, signal_6542, signal_6541, signal_2317}), .clk ( clk ), .r ({Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .c ({signal_6633, signal_6632, signal_6631, signal_2347}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2333 ( .a ({signal_5838, signal_5837, signal_5836, signal_2082}), .b ({signal_6579, signal_6578, signal_6577, signal_2329}), .clk ( clk ), .r ({Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016]}), .c ({signal_6636, signal_6635, signal_6634, signal_2348}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2335 ( .a ({signal_6612, signal_6611, signal_6610, signal_2340}), .b ({signal_6642, signal_6641, signal_6640, signal_2350}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2336 ( .a ({signal_6633, signal_6632, signal_6631, signal_2347}), .b ({signal_6645, signal_6644, signal_6643, signal_2351}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2337 ( .a ({signal_6231, signal_6230, signal_6229, signal_2213}), .b ({signal_6615, signal_6614, signal_6613, signal_2341}), .clk ( clk ), .r ({Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022]}), .c ({signal_6648, signal_6647, signal_6646, signal_2352}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2339 ( .a ({signal_6348, signal_6347, signal_6346, signal_2252}), .b ({signal_6624, signal_6623, signal_6622, signal_2344}), .clk ( clk ), .r ({Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028]}), .c ({signal_6654, signal_6653, signal_6652, signal_2354}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2340 ( .a ({signal_6072, signal_6071, signal_6070, signal_2160}), .b ({signal_6603, signal_6602, signal_6601, signal_2337}), .clk ( clk ), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034]}), .c ({signal_6657, signal_6656, signal_6655, signal_2355}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2341 ( .a ({signal_6159, signal_6158, signal_6157, signal_2189}), .b ({signal_6606, signal_6605, signal_6604, signal_2338}), .clk ( clk ), .r ({Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({signal_6660, signal_6659, signal_6658, signal_2356}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2342 ( .a ({signal_6006, signal_6005, signal_6004, signal_2138}), .b ({signal_6627, signal_6626, signal_6625, signal_2345}), .clk ( clk ), .r ({Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046]}), .c ({signal_6663, signal_6662, signal_6661, signal_2357}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2343 ( .a ({signal_6609, signal_6608, signal_6607, signal_2339}), .b ({signal_6582, signal_6581, signal_6580, signal_2330}), .clk ( clk ), .r ({Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052]}), .c ({signal_6666, signal_6665, signal_6664, signal_2358}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2319 ( .a ({signal_6198, signal_6197, signal_6196, signal_2202}), .b ({signal_6525, signal_6524, signal_6523, signal_2311}), .clk ( clk ), .r ({Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058]}), .c ({signal_6594, signal_6593, signal_6592, signal_2334}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2334 ( .a ({signal_4800, signal_4799, signal_4798, signal_1736}), .b ({signal_6585, signal_6584, signal_6583, signal_2331}), .clk ( clk ), .r ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064]}), .c ({signal_6639, signal_6638, signal_6637, signal_2349}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2338 ( .a ({signal_6306, signal_6305, signal_6304, signal_2238}), .b ({signal_6618, signal_6617, signal_6616, signal_2342}), .clk ( clk ), .r ({Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .c ({signal_6651, signal_6650, signal_6649, signal_2353}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2344 ( .a ({signal_6630, signal_6629, signal_6628, signal_2346}), .b ({signal_6444, signal_6443, signal_6442, signal_2284}), .clk ( clk ), .r ({Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076]}), .c ({signal_6669, signal_6668, signal_6667, signal_2359}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2346 ( .a ({signal_6222, signal_6221, signal_6220, signal_2210}), .b ({signal_6642, signal_6641, signal_6640, signal_2350}), .clk ( clk ), .r ({Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082]}), .c ({signal_6675, signal_6674, signal_6673, signal_2361}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2348 ( .a ({signal_4173, signal_4172, signal_4171, signal_1527}), .b ({signal_6657, signal_6656, signal_6655, signal_2355}), .clk ( clk ), .r ({Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088]}), .c ({signal_6681, signal_6680, signal_6679, signal_2363}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2349 ( .a ({signal_6054, signal_6053, signal_6052, signal_2154}), .b ({signal_6660, signal_6659, signal_6658, signal_2356}), .clk ( clk ), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094]}), .c ({signal_6684, signal_6683, signal_6682, signal_2364}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2350 ( .a ({signal_4491, signal_4490, signal_4489, signal_1633}), .b ({signal_6645, signal_6644, signal_6643, signal_2351}), .clk ( clk ), .r ({Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({signal_6687, signal_6686, signal_6685, signal_2365}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2351 ( .a ({signal_6039, signal_6038, signal_6037, signal_2149}), .b ({signal_6666, signal_6665, signal_6664, signal_2358}), .clk ( clk ), .r ({Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106]}), .c ({signal_6690, signal_6689, signal_6688, signal_2366}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2352 ( .a ({signal_6648, signal_6647, signal_6646, signal_2352}), .b ({signal_6591, signal_6590, signal_6589, signal_2333}), .clk ( clk ), .r ({Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112]}), .c ({signal_6693, signal_6692, signal_6691, signal_2367}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2345 ( .a ({signal_6597, signal_6596, signal_6595, signal_2335}), .b ({signal_6594, signal_6593, signal_6592, signal_2334}), .clk ( clk ), .r ({Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118]}), .c ({signal_6672, signal_6671, signal_6670, signal_2360}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2347 ( .a ({signal_6048, signal_6047, signal_6046, signal_2152}), .b ({signal_6651, signal_6650, signal_6649, signal_2353}), .clk ( clk ), .r ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124]}), .c ({signal_6678, signal_6677, signal_6676, signal_2362}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2353 ( .a ({signal_6654, signal_6653, signal_6652, signal_2354}), .b ({signal_6639, signal_6638, signal_6637, signal_2349}), .clk ( clk ), .r ({Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .c ({signal_6696, signal_6695, signal_6694, signal_2368}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2354 ( .a ({signal_6663, signal_6662, signal_6661, signal_2357}), .b ({signal_6669, signal_6668, signal_6667, signal_2359}), .clk ( clk ), .r ({Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136]}), .c ({signal_6699, signal_6698, signal_6697, signal_2369}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2357 ( .a ({signal_4356, signal_4355, signal_4354, signal_1588}), .b ({signal_6681, signal_6680, signal_6679, signal_2363}), .clk ( clk ), .r ({Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142]}), .c ({signal_6708, signal_6707, signal_6706, signal_2372}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2358 ( .a ({signal_6516, signal_6515, signal_6514, signal_2308}), .b ({signal_6684, signal_6683, signal_6682, signal_2364}), .clk ( clk ), .r ({Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148]}), .c ({signal_6711, signal_6710, signal_6709, signal_2373}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2359 ( .a ({signal_4398, signal_4397, signal_4396, signal_1602}), .b ({signal_6687, signal_6686, signal_6685, signal_2365}), .clk ( clk ), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154]}), .c ({signal_6714, signal_6713, signal_6712, signal_2374}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2360 ( .a ({signal_6363, signal_6362, signal_6361, signal_2257}), .b ({signal_6690, signal_6689, signal_6688, signal_2366}), .clk ( clk ), .r ({Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({signal_6717, signal_6716, signal_6715, signal_2375}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2361 ( .a ({signal_6546, signal_6545, signal_6544, signal_2318}), .b ({signal_6693, signal_6692, signal_6691, signal_2367}), .clk ( clk ), .r ({Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166]}), .c ({signal_6720, signal_6719, signal_6718, signal_2376}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2355 ( .a ({signal_6600, signal_6599, signal_6598, signal_2336}), .b ({signal_6672, signal_6671, signal_6670, signal_2360}), .clk ( clk ), .r ({Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172]}), .c ({signal_6702, signal_6701, signal_6700, signal_2370}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2356 ( .a ({signal_6459, signal_6458, signal_6457, signal_2289}), .b ({signal_6678, signal_6677, signal_6676, signal_2362}), .clk ( clk ), .r ({Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178]}), .c ({signal_6705, signal_6704, signal_6703, signal_2371}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2362 ( .a ({signal_6621, signal_6620, signal_6619, signal_2343}), .b ({signal_6696, signal_6695, signal_6694, signal_2368}), .clk ( clk ), .r ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184]}), .c ({signal_6723, signal_6722, signal_6721, signal_2377}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2363 ( .a ({signal_6387, signal_6386, signal_6385, signal_2265}), .b ({signal_6699, signal_6698, signal_6697, signal_2369}), .clk ( clk ), .r ({Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .c ({signal_6726, signal_6725, signal_6724, signal_2378}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2365 ( .a ({signal_6726, signal_6725, signal_6724, signal_2378}), .b ({signal_6732, signal_6731, signal_6730, signal_26}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2368 ( .a ({signal_4941, signal_4940, signal_4939, signal_1783}), .b ({signal_6708, signal_6707, signal_6706, signal_2372}), .clk ( clk ), .r ({Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196]}), .c ({signal_6741, signal_6740, signal_6739, signal_2381}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2369 ( .a ({signal_4209, signal_4208, signal_4207, signal_1539}), .b ({signal_6714, signal_6713, signal_6712, signal_2374}), .clk ( clk ), .r ({Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202]}), .c ({signal_6744, signal_6743, signal_6742, signal_2382}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2370 ( .a ({signal_6636, signal_6635, signal_6634, signal_2348}), .b ({signal_6717, signal_6716, signal_6715, signal_2375}), .clk ( clk ), .r ({Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208]}), .c ({signal_6747, signal_6746, signal_6745, signal_2383}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2371 ( .a ({signal_6435, signal_6434, signal_6433, signal_2281}), .b ({signal_6720, signal_6719, signal_6718, signal_2376}), .clk ( clk ), .r ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214]}), .c ({signal_6750, signal_6749, signal_6748, signal_2384}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2374 ( .a ({signal_6747, signal_6746, signal_6745, signal_2383}), .b ({signal_6759, signal_6758, signal_6757, signal_28}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2375 ( .a ({signal_6750, signal_6749, signal_6748, signal_2384}), .b ({signal_6762, signal_6761, signal_6760, signal_29}) ) ;

    /* cells in depth 27 */

    /* cells in depth 28 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2364 ( .a ({signal_6510, signal_6509, signal_6508, signal_2306}), .b ({signal_6702, signal_6701, signal_6700, signal_2370}), .clk ( clk ), .r ({Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .c ({signal_6729, signal_6728, signal_6727, signal_2379}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2366 ( .a ({signal_6729, signal_6728, signal_6727, signal_2379}), .b ({signal_6735, signal_6734, signal_6733, signal_23}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2367 ( .a ({signal_6447, signal_6446, signal_6445, signal_2285}), .b ({signal_6705, signal_6704, signal_6703, signal_2371}), .clk ( clk ), .r ({Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226]}), .c ({signal_6738, signal_6737, signal_6736, signal_2380}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2372 ( .a ({signal_6675, signal_6674, signal_6673, signal_2361}), .b ({signal_6723, signal_6722, signal_6721, signal_2377}), .clk ( clk ), .r ({Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232]}), .c ({signal_6753, signal_6752, signal_6751, signal_2385}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2373 ( .a ({signal_6738, signal_6737, signal_6736, signal_2380}), .b ({signal_6756, signal_6755, signal_6754, signal_30}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2376 ( .a ({signal_6753, signal_6752, signal_6751, signal_2385}), .b ({signal_6765, signal_6764, signal_6763, signal_24}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2377 ( .a ({signal_6711, signal_6710, signal_6709, signal_2373}), .b ({signal_6741, signal_6740, signal_6739, signal_2381}), .clk ( clk ), .r ({Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238]}), .c ({signal_6768, signal_6767, signal_6766, signal_2386}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2378 ( .a ({signal_4401, signal_4400, signal_4399, signal_1603}), .b ({signal_6744, signal_6743, signal_6742, signal_2382}), .clk ( clk ), .r ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244]}), .c ({signal_6771, signal_6770, signal_6769, signal_2387}) ) ;

    /* cells in depth 29 */

    /* cells in depth 30 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2379 ( .a ({signal_6588, signal_6587, signal_6586, signal_2332}), .b ({signal_6768, signal_6767, signal_6766, signal_2386}), .clk ( clk ), .r ({Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .c ({signal_6774, signal_6773, signal_6772, signal_2388}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2380 ( .a ({signal_6372, signal_6371, signal_6370, signal_2260}), .b ({signal_6771, signal_6770, signal_6769, signal_2387}), .clk ( clk ), .r ({Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256]}), .c ({signal_6777, signal_6776, signal_6775, signal_2389}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2381 ( .a ({signal_6774, signal_6773, signal_6772, signal_2388}), .b ({signal_6780, signal_6779, signal_6778, signal_25}) ) ;

    /* cells in depth 31 */

    /* cells in depth 32 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2382 ( .a ({signal_6558, signal_6557, signal_6556, signal_2322}), .b ({signal_6777, signal_6776, signal_6775, signal_2389}), .clk ( clk ), .r ({Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262]}), .c ({signal_6783, signal_6782, signal_6781, signal_2390}) ) ;

    /* cells in depth 33 */

    /* cells in depth 34 */
    and_HPC2 #(.security_order(3), .pipeline(0)) cell_2383 ( .a ({signal_6576, signal_6575, signal_6574, signal_2328}), .b ({signal_6783, signal_6782, signal_6781, signal_2390}), .clk ( clk ), .r ({Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268]}), .c ({signal_6786, signal_6785, signal_6784, signal_2391}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) cell_2384 ( .a ({signal_6786, signal_6785, signal_6784, signal_2391}), .b ({signal_6789, signal_6788, signal_6787, signal_27}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) cell_0 ( .clk ( signal_12089 ), .D ({signal_6735, signal_6734, signal_6733, signal_23}), .Q ({SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_1 ( .clk ( signal_12089 ), .D ({signal_6765, signal_6764, signal_6763, signal_24}), .Q ({SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_2 ( .clk ( signal_12089 ), .D ({signal_6780, signal_6779, signal_6778, signal_25}), .Q ({SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_3 ( .clk ( signal_12089 ), .D ({signal_6732, signal_6731, signal_6730, signal_26}), .Q ({SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_4 ( .clk ( signal_12089 ), .D ({signal_6789, signal_6788, signal_6787, signal_27}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_5 ( .clk ( signal_12089 ), .D ({signal_6759, signal_6758, signal_6757, signal_28}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_6 ( .clk ( signal_12089 ), .D ({signal_6762, signal_6761, signal_6760, signal_29}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) cell_7 ( .clk ( signal_12089 ), .D ({signal_6756, signal_6755, signal_6754, signal_30}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
