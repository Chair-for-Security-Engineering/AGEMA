
module SkinnyTop ( clk, rst, Plaintext, Key, Ciphertext, done );
  (* AGEMA = "secure" *) input [63:0] Plaintext;
  (* AGEMA = "secure" *) input [63:0] Key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input rst;

  output [63:0] Ciphertext;
  output done;
  
  wire   StateReg_s_current_state_reg_63__QN,
         StateReg_s_current_state_reg_62__QN,
         StateReg_s_current_state_reg_61__QN,
         StateReg_s_current_state_reg_60__QN,
         StateReg_s_current_state_reg_59__QN,
         StateReg_s_current_state_reg_58__QN,
         StateReg_s_current_state_reg_57__QN,
         StateReg_s_current_state_reg_56__QN,
         StateReg_s_current_state_reg_55__QN,
         StateReg_s_current_state_reg_54__QN,
         StateReg_s_current_state_reg_53__QN,
         StateReg_s_current_state_reg_52__QN,
         StateReg_s_current_state_reg_51__QN,
         StateReg_s_current_state_reg_50__QN,
         StateReg_s_current_state_reg_49__QN,
         StateReg_s_current_state_reg_48__QN,
         StateReg_s_current_state_reg_47__QN,
         StateReg_s_current_state_reg_46__QN,
         StateReg_s_current_state_reg_45__QN,
         StateReg_s_current_state_reg_44__QN,
         StateReg_s_current_state_reg_43__QN,
         StateReg_s_current_state_reg_42__QN,
         StateReg_s_current_state_reg_41__QN,
         StateReg_s_current_state_reg_40__QN,
         StateReg_s_current_state_reg_39__QN,
         StateReg_s_current_state_reg_38__QN,
         StateReg_s_current_state_reg_37__QN,
         StateReg_s_current_state_reg_36__QN,
         StateReg_s_current_state_reg_35__QN,
         StateReg_s_current_state_reg_34__QN,
         StateReg_s_current_state_reg_33__QN,
         StateReg_s_current_state_reg_32__QN,
         StateReg_s_current_state_reg_31__QN,
         StateReg_s_current_state_reg_30__QN,
         StateReg_s_current_state_reg_29__QN,
         StateReg_s_current_state_reg_28__QN,
         StateReg_s_current_state_reg_27__QN,
         StateReg_s_current_state_reg_26__QN,
         StateReg_s_current_state_reg_25__QN,
         StateReg_s_current_state_reg_24__QN,
         StateReg_s_current_state_reg_23__QN,
         StateReg_s_current_state_reg_22__QN,
         StateReg_s_current_state_reg_21__QN,
         StateReg_s_current_state_reg_20__QN,
         StateReg_s_current_state_reg_19__QN,
         StateReg_s_current_state_reg_18__QN,
         StateReg_s_current_state_reg_17__QN,
         StateReg_s_current_state_reg_16__QN,
         StateReg_s_current_state_reg_15__QN,
         StateReg_s_current_state_reg_14__QN,
         StateReg_s_current_state_reg_13__QN,
         StateReg_s_current_state_reg_12__QN,
         StateReg_s_current_state_reg_11__QN,
         StateReg_s_current_state_reg_10__QN,
         StateReg_s_current_state_reg_9__QN,
         StateReg_s_current_state_reg_8__QN,
         StateReg_s_current_state_reg_7__QN,
         StateReg_s_current_state_reg_6__QN,
         StateReg_s_current_state_reg_5__QN,
         StateReg_s_current_state_reg_4__QN,
         StateReg_s_current_state_reg_3__QN,
         StateReg_s_current_state_reg_2__QN,
         StateReg_s_current_state_reg_1__QN,
         StateReg_s_current_state_reg_0__QN, SubCellInst_SboxInst_0_n3,
         SubCellInst_SboxInst_0_YY_0_, SubCellInst_SboxInst_0_YY_1_,
         SubCellInst_SboxInst_0_L3, SubCellInst_SboxInst_0_YY_3,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_0_T3,
         SubCellInst_SboxInst_0_Q7, SubCellInst_SboxInst_0_L1,
         SubCellInst_SboxInst_0_Q6, SubCellInst_SboxInst_0_L0,
         SubCellInst_SboxInst_0_T2, SubCellInst_SboxInst_0_Q4,
         SubCellInst_SboxInst_0_T1, SubCellInst_SboxInst_0_Q2,
         SubCellInst_SboxInst_0_T0, SubCellInst_SboxInst_0_Q1,
         SubCellInst_SboxInst_0_Q0, SubCellInst_SboxInst_0_XX_1_,
         SubCellInst_SboxInst_0_XX_2_, SubCellInst_SboxInst_1_n3,
         SubCellInst_SboxInst_1_YY_0_, SubCellInst_SboxInst_1_YY_1_,
         SubCellInst_SboxInst_1_L3, SubCellInst_SboxInst_1_YY_3,
         SubCellInst_SboxInst_1_L2, SubCellInst_SboxInst_1_T3,
         SubCellInst_SboxInst_1_Q7, SubCellInst_SboxInst_1_L1,
         SubCellInst_SboxInst_1_Q6, SubCellInst_SboxInst_1_L0,
         SubCellInst_SboxInst_1_T2, SubCellInst_SboxInst_1_Q4,
         SubCellInst_SboxInst_1_T1, SubCellInst_SboxInst_1_Q2,
         SubCellInst_SboxInst_1_T0, SubCellInst_SboxInst_1_Q1,
         SubCellInst_SboxInst_1_Q0, SubCellInst_SboxInst_1_XX_1_,
         SubCellInst_SboxInst_1_XX_2_, SubCellInst_SboxInst_2_n3,
         SubCellInst_SboxInst_2_YY_0_, SubCellInst_SboxInst_2_YY_1_,
         SubCellInst_SboxInst_2_L3, SubCellInst_SboxInst_2_YY_3,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_2_T3,
         SubCellInst_SboxInst_2_Q7, SubCellInst_SboxInst_2_L1,
         SubCellInst_SboxInst_2_Q6, SubCellInst_SboxInst_2_L0,
         SubCellInst_SboxInst_2_T2, SubCellInst_SboxInst_2_Q4,
         SubCellInst_SboxInst_2_T1, SubCellInst_SboxInst_2_Q2,
         SubCellInst_SboxInst_2_T0, SubCellInst_SboxInst_2_Q1,
         SubCellInst_SboxInst_2_Q0, SubCellInst_SboxInst_2_XX_1_,
         SubCellInst_SboxInst_2_XX_2_, SubCellInst_SboxInst_3_n3,
         SubCellInst_SboxInst_3_YY_0_, SubCellInst_SboxInst_3_YY_1_,
         SubCellInst_SboxInst_3_L3, SubCellInst_SboxInst_3_YY_3,
         SubCellInst_SboxInst_3_L2, SubCellInst_SboxInst_3_T3,
         SubCellInst_SboxInst_3_Q7, SubCellInst_SboxInst_3_L1,
         SubCellInst_SboxInst_3_Q6, SubCellInst_SboxInst_3_L0,
         SubCellInst_SboxInst_3_T2, SubCellInst_SboxInst_3_Q4,
         SubCellInst_SboxInst_3_T1, SubCellInst_SboxInst_3_Q2,
         SubCellInst_SboxInst_3_T0, SubCellInst_SboxInst_3_Q1,
         SubCellInst_SboxInst_3_Q0, SubCellInst_SboxInst_3_XX_1_,
         SubCellInst_SboxInst_3_XX_2_, SubCellInst_SboxInst_4_n3,
         SubCellInst_SboxInst_4_YY_0_, SubCellInst_SboxInst_4_YY_1_,
         SubCellInst_SboxInst_4_L3, SubCellInst_SboxInst_4_YY_3,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_4_T3,
         SubCellInst_SboxInst_4_Q7, SubCellInst_SboxInst_4_L1,
         SubCellInst_SboxInst_4_Q6, SubCellInst_SboxInst_4_L0,
         SubCellInst_SboxInst_4_T2, SubCellInst_SboxInst_4_Q4,
         SubCellInst_SboxInst_4_T1, SubCellInst_SboxInst_4_Q2,
         SubCellInst_SboxInst_4_T0, SubCellInst_SboxInst_4_Q1,
         SubCellInst_SboxInst_4_Q0, SubCellInst_SboxInst_4_XX_1_,
         SubCellInst_SboxInst_4_XX_2_, SubCellInst_SboxInst_5_n3,
         SubCellInst_SboxInst_5_YY_0_, SubCellInst_SboxInst_5_YY_1_,
         SubCellInst_SboxInst_5_L3, SubCellInst_SboxInst_5_YY_3,
         SubCellInst_SboxInst_5_L2, SubCellInst_SboxInst_5_T3,
         SubCellInst_SboxInst_5_Q7, SubCellInst_SboxInst_5_L1,
         SubCellInst_SboxInst_5_Q6, SubCellInst_SboxInst_5_L0,
         SubCellInst_SboxInst_5_T2, SubCellInst_SboxInst_5_Q4,
         SubCellInst_SboxInst_5_T1, SubCellInst_SboxInst_5_Q2,
         SubCellInst_SboxInst_5_T0, SubCellInst_SboxInst_5_Q1,
         SubCellInst_SboxInst_5_Q0, SubCellInst_SboxInst_5_XX_1_,
         SubCellInst_SboxInst_5_XX_2_, SubCellInst_SboxInst_6_n3,
         SubCellInst_SboxInst_6_YY_0_, SubCellInst_SboxInst_6_YY_1_,
         SubCellInst_SboxInst_6_L3, SubCellInst_SboxInst_6_YY_3,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_6_T3,
         SubCellInst_SboxInst_6_Q7, SubCellInst_SboxInst_6_L1,
         SubCellInst_SboxInst_6_Q6, SubCellInst_SboxInst_6_L0,
         SubCellInst_SboxInst_6_T2, SubCellInst_SboxInst_6_Q4,
         SubCellInst_SboxInst_6_T1, SubCellInst_SboxInst_6_Q2,
         SubCellInst_SboxInst_6_T0, SubCellInst_SboxInst_6_Q1,
         SubCellInst_SboxInst_6_Q0, SubCellInst_SboxInst_6_XX_1_,
         SubCellInst_SboxInst_6_XX_2_, SubCellInst_SboxInst_7_n3,
         SubCellInst_SboxInst_7_YY_0_, SubCellInst_SboxInst_7_YY_1_,
         SubCellInst_SboxInst_7_L3, SubCellInst_SboxInst_7_YY_3,
         SubCellInst_SboxInst_7_L2, SubCellInst_SboxInst_7_T3,
         SubCellInst_SboxInst_7_Q7, SubCellInst_SboxInst_7_L1,
         SubCellInst_SboxInst_7_Q6, SubCellInst_SboxInst_7_L0,
         SubCellInst_SboxInst_7_T2, SubCellInst_SboxInst_7_Q4,
         SubCellInst_SboxInst_7_T1, SubCellInst_SboxInst_7_Q2,
         SubCellInst_SboxInst_7_T0, SubCellInst_SboxInst_7_Q1,
         SubCellInst_SboxInst_7_Q0, SubCellInst_SboxInst_7_XX_1_,
         SubCellInst_SboxInst_7_XX_2_, SubCellInst_SboxInst_8_n3,
         SubCellInst_SboxInst_8_YY_0_, SubCellInst_SboxInst_8_YY_1_,
         SubCellInst_SboxInst_8_L3, SubCellInst_SboxInst_8_YY_3,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_8_T3,
         SubCellInst_SboxInst_8_Q7, SubCellInst_SboxInst_8_L1,
         SubCellInst_SboxInst_8_Q6, SubCellInst_SboxInst_8_L0,
         SubCellInst_SboxInst_8_T2, SubCellInst_SboxInst_8_Q4,
         SubCellInst_SboxInst_8_T1, SubCellInst_SboxInst_8_Q2,
         SubCellInst_SboxInst_8_T0, SubCellInst_SboxInst_8_Q1,
         SubCellInst_SboxInst_8_Q0, SubCellInst_SboxInst_8_XX_1_,
         SubCellInst_SboxInst_8_XX_2_, SubCellInst_SboxInst_9_n3,
         SubCellInst_SboxInst_9_YY_0_, SubCellInst_SboxInst_9_YY_1_,
         SubCellInst_SboxInst_9_L3, SubCellInst_SboxInst_9_YY_3,
         SubCellInst_SboxInst_9_L2, SubCellInst_SboxInst_9_T3,
         SubCellInst_SboxInst_9_Q7, SubCellInst_SboxInst_9_L1,
         SubCellInst_SboxInst_9_Q6, SubCellInst_SboxInst_9_L0,
         SubCellInst_SboxInst_9_T2, SubCellInst_SboxInst_9_Q4,
         SubCellInst_SboxInst_9_T1, SubCellInst_SboxInst_9_Q2,
         SubCellInst_SboxInst_9_T0, SubCellInst_SboxInst_9_Q1,
         SubCellInst_SboxInst_9_Q0, SubCellInst_SboxInst_9_XX_1_,
         SubCellInst_SboxInst_9_XX_2_, SubCellInst_SboxInst_10_n3,
         SubCellInst_SboxInst_10_YY_0_, SubCellInst_SboxInst_10_YY_1_,
         SubCellInst_SboxInst_10_L3, SubCellInst_SboxInst_10_YY_3,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_10_T3,
         SubCellInst_SboxInst_10_Q7, SubCellInst_SboxInst_10_L1,
         SubCellInst_SboxInst_10_Q6, SubCellInst_SboxInst_10_L0,
         SubCellInst_SboxInst_10_T2, SubCellInst_SboxInst_10_Q4,
         SubCellInst_SboxInst_10_T1, SubCellInst_SboxInst_10_Q2,
         SubCellInst_SboxInst_10_T0, SubCellInst_SboxInst_10_Q1,
         SubCellInst_SboxInst_10_Q0, SubCellInst_SboxInst_10_XX_1_,
         SubCellInst_SboxInst_10_XX_2_, SubCellInst_SboxInst_11_n3,
         SubCellInst_SboxInst_11_YY_0_, SubCellInst_SboxInst_11_YY_1_,
         SubCellInst_SboxInst_11_L3, SubCellInst_SboxInst_11_YY_3,
         SubCellInst_SboxInst_11_L2, SubCellInst_SboxInst_11_T3,
         SubCellInst_SboxInst_11_Q7, SubCellInst_SboxInst_11_L1,
         SubCellInst_SboxInst_11_Q6, SubCellInst_SboxInst_11_L0,
         SubCellInst_SboxInst_11_T2, SubCellInst_SboxInst_11_Q4,
         SubCellInst_SboxInst_11_T1, SubCellInst_SboxInst_11_Q2,
         SubCellInst_SboxInst_11_T0, SubCellInst_SboxInst_11_Q1,
         SubCellInst_SboxInst_11_Q0, SubCellInst_SboxInst_11_XX_1_,
         SubCellInst_SboxInst_11_XX_2_, SubCellInst_SboxInst_12_n3,
         SubCellInst_SboxInst_12_YY_0_, SubCellInst_SboxInst_12_YY_1_,
         SubCellInst_SboxInst_12_L3, SubCellInst_SboxInst_12_YY_3,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_12_T3,
         SubCellInst_SboxInst_12_Q7, SubCellInst_SboxInst_12_L1,
         SubCellInst_SboxInst_12_Q6, SubCellInst_SboxInst_12_L0,
         SubCellInst_SboxInst_12_T2, SubCellInst_SboxInst_12_Q4,
         SubCellInst_SboxInst_12_T1, SubCellInst_SboxInst_12_Q2,
         SubCellInst_SboxInst_12_T0, SubCellInst_SboxInst_12_Q1,
         SubCellInst_SboxInst_12_Q0, SubCellInst_SboxInst_12_XX_1_,
         SubCellInst_SboxInst_12_XX_2_, SubCellInst_SboxInst_13_n3,
         SubCellInst_SboxInst_13_YY_0_, SubCellInst_SboxInst_13_YY_1_,
         SubCellInst_SboxInst_13_L3, SubCellInst_SboxInst_13_YY_3,
         SubCellInst_SboxInst_13_L2, SubCellInst_SboxInst_13_T3,
         SubCellInst_SboxInst_13_Q7, SubCellInst_SboxInst_13_L1,
         SubCellInst_SboxInst_13_Q6, SubCellInst_SboxInst_13_L0,
         SubCellInst_SboxInst_13_T2, SubCellInst_SboxInst_13_Q4,
         SubCellInst_SboxInst_13_T1, SubCellInst_SboxInst_13_Q2,
         SubCellInst_SboxInst_13_T0, SubCellInst_SboxInst_13_Q1,
         SubCellInst_SboxInst_13_Q0, SubCellInst_SboxInst_13_XX_1_,
         SubCellInst_SboxInst_13_XX_2_, SubCellInst_SboxInst_14_n3,
         SubCellInst_SboxInst_14_YY_0_, SubCellInst_SboxInst_14_YY_1_,
         SubCellInst_SboxInst_14_L3, SubCellInst_SboxInst_14_YY_3,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_14_T3,
         SubCellInst_SboxInst_14_Q7, SubCellInst_SboxInst_14_L1,
         SubCellInst_SboxInst_14_Q6, SubCellInst_SboxInst_14_L0,
         SubCellInst_SboxInst_14_T2, SubCellInst_SboxInst_14_Q4,
         SubCellInst_SboxInst_14_T1, SubCellInst_SboxInst_14_Q2,
         SubCellInst_SboxInst_14_T0, SubCellInst_SboxInst_14_Q1,
         SubCellInst_SboxInst_14_Q0, SubCellInst_SboxInst_14_XX_1_,
         SubCellInst_SboxInst_14_XX_2_, SubCellInst_SboxInst_15_n3,
         SubCellInst_SboxInst_15_YY_0_, SubCellInst_SboxInst_15_YY_1_,
         SubCellInst_SboxInst_15_L3, SubCellInst_SboxInst_15_YY_3,
         SubCellInst_SboxInst_15_L2, SubCellInst_SboxInst_15_T3,
         SubCellInst_SboxInst_15_Q7, SubCellInst_SboxInst_15_L1,
         SubCellInst_SboxInst_15_Q6, SubCellInst_SboxInst_15_L0,
         SubCellInst_SboxInst_15_T2, SubCellInst_SboxInst_15_Q4,
         SubCellInst_SboxInst_15_T1, SubCellInst_SboxInst_15_Q2,
         SubCellInst_SboxInst_15_T0, SubCellInst_SboxInst_15_Q1,
         SubCellInst_SboxInst_15_Q0, SubCellInst_SboxInst_15_XX_1_,
         SubCellInst_SboxInst_15_XX_2_, AddConstXOR_AddConstXOR_XORInst_0_0_n1,
         AddConstXOR_AddConstXOR_XORInst_0_1_n1,
         AddConstXOR_AddConstXOR_XORInst_0_2_n1,
         AddConstXOR_AddConstXOR_XORInst_0_3_n1,
         AddConstXOR_AddConstXOR_XORInst_1_0_n1,
         AddConstXOR_AddConstXOR_XORInst_1_1_n1,
         AddConstXOR_AddConstXOR_XORInst_1_2_n1,
         AddConstXOR_AddConstXOR_XORInst_1_3_n1,
         AddRoundTweakeyXOR_XORInst_0_0_n1, AddRoundTweakeyXOR_XORInst_0_1_n1,
         AddRoundTweakeyXOR_XORInst_0_2_n1, AddRoundTweakeyXOR_XORInst_0_3_n1,
         AddRoundTweakeyXOR_XORInst_1_0_n1, AddRoundTweakeyXOR_XORInst_1_1_n1,
         AddRoundTweakeyXOR_XORInst_1_2_n1, AddRoundTweakeyXOR_XORInst_1_3_n1,
         AddRoundTweakeyXOR_XORInst_2_0_n1, AddRoundTweakeyXOR_XORInst_2_1_n1,
         AddRoundTweakeyXOR_XORInst_2_2_n1, AddRoundTweakeyXOR_XORInst_2_3_n1,
         AddRoundTweakeyXOR_XORInst_3_0_n1, AddRoundTweakeyXOR_XORInst_3_1_n1,
         AddRoundTweakeyXOR_XORInst_3_2_n1, AddRoundTweakeyXOR_XORInst_3_3_n1,
         AddRoundTweakeyXOR_XORInst_4_0_n1, AddRoundTweakeyXOR_XORInst_4_1_n1,
         AddRoundTweakeyXOR_XORInst_4_2_n1, AddRoundTweakeyXOR_XORInst_4_3_n1,
         AddRoundTweakeyXOR_XORInst_5_0_n1, AddRoundTweakeyXOR_XORInst_5_1_n1,
         AddRoundTweakeyXOR_XORInst_5_2_n1, AddRoundTweakeyXOR_XORInst_5_3_n1,
         AddRoundTweakeyXOR_XORInst_6_0_n1, AddRoundTweakeyXOR_XORInst_6_1_n1,
         AddRoundTweakeyXOR_XORInst_6_2_n1, AddRoundTweakeyXOR_XORInst_6_3_n1,
         AddRoundTweakeyXOR_XORInst_7_0_n1, AddRoundTweakeyXOR_XORInst_7_1_n1,
         AddRoundTweakeyXOR_XORInst_7_2_n1, AddRoundTweakeyXOR_XORInst_7_3_n1,
         MCInst_MCR0_XORInst_0_0_n2, MCInst_MCR0_XORInst_0_0_n1,
         MCInst_MCR0_XORInst_0_1_n2, MCInst_MCR0_XORInst_0_1_n1,
         MCInst_MCR0_XORInst_0_2_n2, MCInst_MCR0_XORInst_0_2_n1,
         MCInst_MCR0_XORInst_0_3_n2, MCInst_MCR0_XORInst_0_3_n1,
         MCInst_MCR0_XORInst_1_0_n2, MCInst_MCR0_XORInst_1_0_n1,
         MCInst_MCR0_XORInst_1_1_n2, MCInst_MCR0_XORInst_1_1_n1,
         MCInst_MCR0_XORInst_1_2_n2, MCInst_MCR0_XORInst_1_2_n1,
         MCInst_MCR0_XORInst_1_3_n2, MCInst_MCR0_XORInst_1_3_n1,
         MCInst_MCR0_XORInst_2_0_n2, MCInst_MCR0_XORInst_2_0_n1,
         MCInst_MCR0_XORInst_2_1_n2, MCInst_MCR0_XORInst_2_1_n1,
         MCInst_MCR0_XORInst_2_2_n2, MCInst_MCR0_XORInst_2_2_n1,
         MCInst_MCR0_XORInst_2_3_n2, MCInst_MCR0_XORInst_2_3_n1,
         MCInst_MCR0_XORInst_3_0_n2, MCInst_MCR0_XORInst_3_0_n1,
         MCInst_MCR0_XORInst_3_1_n2, MCInst_MCR0_XORInst_3_1_n1,
         MCInst_MCR0_XORInst_3_2_n2, MCInst_MCR0_XORInst_3_2_n1,
         MCInst_MCR0_XORInst_3_3_n2, MCInst_MCR0_XORInst_3_3_n1,
         MCInst_MCR2_XORInst_0_0_n1, MCInst_MCR2_XORInst_0_1_n1,
         MCInst_MCR2_XORInst_0_2_n1, MCInst_MCR2_XORInst_0_3_n1,
         MCInst_MCR2_XORInst_1_0_n1, MCInst_MCR2_XORInst_1_1_n1,
         MCInst_MCR2_XORInst_1_2_n1, MCInst_MCR2_XORInst_1_3_n1,
         MCInst_MCR2_XORInst_2_0_n1, MCInst_MCR2_XORInst_2_1_n1,
         MCInst_MCR2_XORInst_2_2_n1, MCInst_MCR2_XORInst_2_3_n1,
         MCInst_MCR2_XORInst_3_0_n1, MCInst_MCR2_XORInst_3_1_n1,
         MCInst_MCR2_XORInst_3_2_n1, MCInst_MCR2_XORInst_3_3_n1,
         MCInst_MCR3_XORInst_0_0_n1, MCInst_MCR3_XORInst_0_1_n1,
         MCInst_MCR3_XORInst_0_2_n1, MCInst_MCR3_XORInst_0_3_n1,
         MCInst_MCR3_XORInst_1_0_n1, MCInst_MCR3_XORInst_1_1_n1,
         MCInst_MCR3_XORInst_1_2_n1, MCInst_MCR3_XORInst_1_3_n1,
         MCInst_MCR3_XORInst_2_0_n1, MCInst_MCR3_XORInst_2_1_n1,
         MCInst_MCR3_XORInst_2_2_n1, MCInst_MCR3_XORInst_2_3_n1,
         MCInst_MCR3_XORInst_3_0_n1, MCInst_MCR3_XORInst_3_1_n1,
         MCInst_MCR3_XORInst_3_2_n1, MCInst_MCR3_XORInst_3_3_n1,
         TweakeyGeneration_StateReg_s_current_state_reg_63__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_62__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_61__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_60__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_59__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_58__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_57__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_56__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_55__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_54__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_53__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_52__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_51__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_50__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_49__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_48__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_47__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_46__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_45__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_44__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_43__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_42__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_41__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_40__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_39__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_38__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_37__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_36__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_35__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_34__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_33__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_32__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_31__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_30__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_29__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_28__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_27__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_26__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_25__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_24__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_23__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_22__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_21__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_20__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_19__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_18__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_17__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_16__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_15__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_14__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_13__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_12__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_11__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_10__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_9__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_8__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_7__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_6__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_5__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_4__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_3__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_2__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_1__QN,
         TweakeyGeneration_StateReg_s_current_state_reg_0__QN,
         FSMReg_s_current_state_reg_5__QN, FSMReg_s_current_state_reg_4__QN,
         FSMReg_s_current_state_reg_3__QN, FSMReg_s_current_state_reg_2__QN,
         FSMReg_s_current_state_reg_1__QN, FSMReg_s_current_state_reg_0__QN,
         FSMUpdateInst_StateUpdateInst_0_n4,
         FSMUpdateInst_StateUpdateInst_0_n3,
         FSMUpdateInst_StateUpdateInst_0_n2,
         FSMUpdateInst_StateUpdateInst_0_n1,
         FSMUpdateInst_StateUpdateInst_2_n4,
         FSMUpdateInst_StateUpdateInst_2_n3,
         FSMUpdateInst_StateUpdateInst_2_n2,
         FSMUpdateInst_StateUpdateInst_2_n1,
         FSMUpdateInst_StateUpdateInst_5_n4,
         FSMUpdateInst_StateUpdateInst_5_n3,
         FSMUpdateInst_StateUpdateInst_5_n2,
         FSMUpdateInst_StateUpdateInst_5_n1, FSMSignalsInst_doneInst_n5,
         FSMSignalsInst_doneInst_n4, FSMSignalsInst_doneInst_n3,
         FSMSignalsInst_doneInst_n2, FSMSignalsInst_doneInst_n1;
  wire   [63:0] MCOutput;
  wire   [63:0] StateRegInput;
  wire   [63:29] SubCellOutput;
  wire   [5:1] FSM;
  wire   [63:32] AddRoundConstantOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [5:0] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;

  MUX2_X1 PlaintextMUX_MUXInst_0_U1 ( .A(MCOutput[0]), .B(Plaintext[0]), .S(
        rst), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1 ( .A(MCOutput[1]), .B(Plaintext[1]), .S(
        rst), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1 ( .A(MCOutput[2]), .B(Plaintext[2]), .S(
        rst), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1 ( .A(MCOutput[3]), .B(Plaintext[3]), .S(
        rst), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1 ( .A(MCOutput[4]), .B(Plaintext[4]), .S(
        rst), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1 ( .A(MCOutput[5]), .B(Plaintext[5]), .S(
        rst), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1 ( .A(MCOutput[6]), .B(Plaintext[6]), .S(
        rst), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1 ( .A(MCOutput[7]), .B(Plaintext[7]), .S(
        rst), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1 ( .A(MCOutput[8]), .B(Plaintext[8]), .S(
        rst), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1 ( .A(MCOutput[9]), .B(Plaintext[9]), .S(
        rst), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1 ( .A(MCOutput[10]), .B(Plaintext[10]), 
        .S(rst), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1 ( .A(MCOutput[11]), .B(Plaintext[11]), 
        .S(rst), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1 ( .A(MCOutput[12]), .B(Plaintext[12]), 
        .S(rst), .Z(StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1 ( .A(MCOutput[13]), .B(Plaintext[13]), 
        .S(rst), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1 ( .A(MCOutput[14]), .B(Plaintext[14]), 
        .S(rst), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1 ( .A(MCOutput[15]), .B(Plaintext[15]), 
        .S(rst), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1 ( .A(MCOutput[16]), .B(Plaintext[16]), 
        .S(rst), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1 ( .A(MCOutput[17]), .B(Plaintext[17]), 
        .S(rst), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1 ( .A(MCOutput[18]), .B(Plaintext[18]), 
        .S(rst), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1 ( .A(MCOutput[19]), .B(Plaintext[19]), 
        .S(rst), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1 ( .A(MCOutput[20]), .B(Plaintext[20]), 
        .S(rst), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1 ( .A(MCOutput[21]), .B(Plaintext[21]), 
        .S(rst), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1 ( .A(MCOutput[22]), .B(Plaintext[22]), 
        .S(rst), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1 ( .A(MCOutput[23]), .B(Plaintext[23]), 
        .S(rst), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1 ( .A(MCOutput[24]), .B(Plaintext[24]), 
        .S(rst), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1 ( .A(MCOutput[25]), .B(Plaintext[25]), 
        .S(rst), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1 ( .A(MCOutput[26]), .B(Plaintext[26]), 
        .S(rst), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1 ( .A(MCOutput[27]), .B(Plaintext[27]), 
        .S(rst), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1 ( .A(MCOutput[28]), .B(Plaintext[28]), 
        .S(rst), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1 ( .A(MCOutput[29]), .B(Plaintext[29]), 
        .S(rst), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1 ( .A(MCOutput[30]), .B(Plaintext[30]), 
        .S(rst), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1 ( .A(MCOutput[31]), .B(Plaintext[31]), 
        .S(rst), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1 ( .A(MCOutput[32]), .B(Plaintext[32]), 
        .S(rst), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1 ( .A(MCOutput[33]), .B(Plaintext[33]), 
        .S(rst), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1 ( .A(MCOutput[34]), .B(Plaintext[34]), 
        .S(rst), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1 ( .A(MCOutput[35]), .B(Plaintext[35]), 
        .S(rst), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1 ( .A(MCOutput[36]), .B(Plaintext[36]), 
        .S(rst), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1 ( .A(MCOutput[37]), .B(Plaintext[37]), 
        .S(rst), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1 ( .A(MCOutput[38]), .B(Plaintext[38]), 
        .S(rst), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1 ( .A(MCOutput[39]), .B(Plaintext[39]), 
        .S(rst), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1 ( .A(MCOutput[40]), .B(Plaintext[40]), 
        .S(rst), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1 ( .A(MCOutput[41]), .B(Plaintext[41]), 
        .S(rst), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1 ( .A(MCOutput[42]), .B(Plaintext[42]), 
        .S(rst), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1 ( .A(MCOutput[43]), .B(Plaintext[43]), 
        .S(rst), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1 ( .A(MCOutput[44]), .B(Plaintext[44]), 
        .S(rst), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1 ( .A(MCOutput[45]), .B(Plaintext[45]), 
        .S(rst), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1 ( .A(MCOutput[46]), .B(Plaintext[46]), 
        .S(rst), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1 ( .A(MCOutput[47]), .B(Plaintext[47]), 
        .S(rst), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1 ( .A(MCOutput[48]), .B(Plaintext[48]), 
        .S(rst), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1 ( .A(MCOutput[49]), .B(Plaintext[49]), 
        .S(rst), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1 ( .A(MCOutput[50]), .B(Plaintext[50]), 
        .S(rst), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1 ( .A(MCOutput[51]), .B(Plaintext[51]), 
        .S(rst), .Z(StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1 ( .A(MCOutput[52]), .B(Plaintext[52]), 
        .S(rst), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1 ( .A(MCOutput[53]), .B(Plaintext[53]), 
        .S(rst), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1 ( .A(MCOutput[54]), .B(Plaintext[54]), 
        .S(rst), .Z(StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1 ( .A(MCOutput[55]), .B(Plaintext[55]), 
        .S(rst), .Z(StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1 ( .A(MCOutput[56]), .B(Plaintext[56]), 
        .S(rst), .Z(StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1 ( .A(MCOutput[57]), .B(Plaintext[57]), 
        .S(rst), .Z(StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1 ( .A(MCOutput[58]), .B(Plaintext[58]), 
        .S(rst), .Z(StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1 ( .A(MCOutput[59]), .B(Plaintext[59]), 
        .S(rst), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1 ( .A(MCOutput[60]), .B(Plaintext[60]), 
        .S(rst), .Z(StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1 ( .A(MCOutput[61]), .B(Plaintext[61]), 
        .S(rst), .Z(StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1 ( .A(MCOutput[62]), .B(Plaintext[62]), 
        .S(rst), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1 ( .A(MCOutput[63]), .B(Plaintext[63]), 
        .S(rst), .Z(StateRegInput[63]) );
  INV_X1 StateReg_s_current_state_reg_63__U1 ( .A(Ciphertext[63]), .ZN(
        StateReg_s_current_state_reg_63__QN) );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF ( .D(StateRegInput[63]), .CK(
        clk), .Q(Ciphertext[63]), .QN() );
  INV_X1 StateReg_s_current_state_reg_62__U1 ( .A(Ciphertext[62]), .ZN(
        StateReg_s_current_state_reg_62__QN) );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF ( .D(StateRegInput[62]), .CK(
        clk), .Q(Ciphertext[62]), .QN() );
  INV_X1 StateReg_s_current_state_reg_61__U1 ( .A(Ciphertext[61]), .ZN(
        StateReg_s_current_state_reg_61__QN) );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF ( .D(StateRegInput[61]), .CK(
        clk), .Q(Ciphertext[61]), .QN() );
  INV_X1 StateReg_s_current_state_reg_60__U1 ( .A(Ciphertext[60]), .ZN(
        StateReg_s_current_state_reg_60__QN) );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF ( .D(StateRegInput[60]), .CK(
        clk), .Q(Ciphertext[60]), .QN() );
  INV_X1 StateReg_s_current_state_reg_59__U1 ( .A(Ciphertext[59]), .ZN(
        StateReg_s_current_state_reg_59__QN) );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF ( .D(StateRegInput[59]), .CK(
        clk), .Q(Ciphertext[59]), .QN() );
  INV_X1 StateReg_s_current_state_reg_58__U1 ( .A(Ciphertext[58]), .ZN(
        StateReg_s_current_state_reg_58__QN) );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF ( .D(StateRegInput[58]), .CK(
        clk), .Q(Ciphertext[58]), .QN() );
  INV_X1 StateReg_s_current_state_reg_57__U1 ( .A(Ciphertext[57]), .ZN(
        StateReg_s_current_state_reg_57__QN) );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF ( .D(StateRegInput[57]), .CK(
        clk), .Q(Ciphertext[57]), .QN() );
  INV_X1 StateReg_s_current_state_reg_56__U1 ( .A(Ciphertext[56]), .ZN(
        StateReg_s_current_state_reg_56__QN) );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF ( .D(StateRegInput[56]), .CK(
        clk), .Q(Ciphertext[56]), .QN() );
  INV_X1 StateReg_s_current_state_reg_55__U1 ( .A(Ciphertext[55]), .ZN(
        StateReg_s_current_state_reg_55__QN) );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF ( .D(StateRegInput[55]), .CK(
        clk), .Q(Ciphertext[55]), .QN() );
  INV_X1 StateReg_s_current_state_reg_54__U1 ( .A(Ciphertext[54]), .ZN(
        StateReg_s_current_state_reg_54__QN) );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF ( .D(StateRegInput[54]), .CK(
        clk), .Q(Ciphertext[54]), .QN() );
  INV_X1 StateReg_s_current_state_reg_53__U1 ( .A(Ciphertext[53]), .ZN(
        StateReg_s_current_state_reg_53__QN) );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF ( .D(StateRegInput[53]), .CK(
        clk), .Q(Ciphertext[53]), .QN() );
  INV_X1 StateReg_s_current_state_reg_52__U1 ( .A(Ciphertext[52]), .ZN(
        StateReg_s_current_state_reg_52__QN) );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF ( .D(StateRegInput[52]), .CK(
        clk), .Q(Ciphertext[52]), .QN() );
  INV_X1 StateReg_s_current_state_reg_51__U1 ( .A(Ciphertext[51]), .ZN(
        StateReg_s_current_state_reg_51__QN) );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF ( .D(StateRegInput[51]), .CK(
        clk), .Q(Ciphertext[51]), .QN() );
  INV_X1 StateReg_s_current_state_reg_50__U1 ( .A(Ciphertext[50]), .ZN(
        StateReg_s_current_state_reg_50__QN) );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF ( .D(StateRegInput[50]), .CK(
        clk), .Q(Ciphertext[50]), .QN() );
  INV_X1 StateReg_s_current_state_reg_49__U1 ( .A(Ciphertext[49]), .ZN(
        StateReg_s_current_state_reg_49__QN) );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF ( .D(StateRegInput[49]), .CK(
        clk), .Q(Ciphertext[49]), .QN() );
  INV_X1 StateReg_s_current_state_reg_48__U1 ( .A(Ciphertext[48]), .ZN(
        StateReg_s_current_state_reg_48__QN) );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF ( .D(StateRegInput[48]), .CK(
        clk), .Q(Ciphertext[48]), .QN() );
  INV_X1 StateReg_s_current_state_reg_47__U1 ( .A(Ciphertext[47]), .ZN(
        StateReg_s_current_state_reg_47__QN) );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF ( .D(StateRegInput[47]), .CK(
        clk), .Q(Ciphertext[47]), .QN() );
  INV_X1 StateReg_s_current_state_reg_46__U1 ( .A(Ciphertext[46]), .ZN(
        StateReg_s_current_state_reg_46__QN) );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF ( .D(StateRegInput[46]), .CK(
        clk), .Q(Ciphertext[46]), .QN() );
  INV_X1 StateReg_s_current_state_reg_45__U1 ( .A(Ciphertext[45]), .ZN(
        StateReg_s_current_state_reg_45__QN) );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF ( .D(StateRegInput[45]), .CK(
        clk), .Q(Ciphertext[45]), .QN() );
  INV_X1 StateReg_s_current_state_reg_44__U1 ( .A(Ciphertext[44]), .ZN(
        StateReg_s_current_state_reg_44__QN) );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF ( .D(StateRegInput[44]), .CK(
        clk), .Q(Ciphertext[44]), .QN() );
  INV_X1 StateReg_s_current_state_reg_43__U1 ( .A(Ciphertext[43]), .ZN(
        StateReg_s_current_state_reg_43__QN) );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF ( .D(StateRegInput[43]), .CK(
        clk), .Q(Ciphertext[43]), .QN() );
  INV_X1 StateReg_s_current_state_reg_42__U1 ( .A(Ciphertext[42]), .ZN(
        StateReg_s_current_state_reg_42__QN) );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF ( .D(StateRegInput[42]), .CK(
        clk), .Q(Ciphertext[42]), .QN() );
  INV_X1 StateReg_s_current_state_reg_41__U1 ( .A(Ciphertext[41]), .ZN(
        StateReg_s_current_state_reg_41__QN) );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF ( .D(StateRegInput[41]), .CK(
        clk), .Q(Ciphertext[41]), .QN() );
  INV_X1 StateReg_s_current_state_reg_40__U1 ( .A(Ciphertext[40]), .ZN(
        StateReg_s_current_state_reg_40__QN) );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF ( .D(StateRegInput[40]), .CK(
        clk), .Q(Ciphertext[40]), .QN() );
  INV_X1 StateReg_s_current_state_reg_39__U1 ( .A(Ciphertext[39]), .ZN(
        StateReg_s_current_state_reg_39__QN) );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF ( .D(StateRegInput[39]), .CK(
        clk), .Q(Ciphertext[39]), .QN() );
  INV_X1 StateReg_s_current_state_reg_38__U1 ( .A(Ciphertext[38]), .ZN(
        StateReg_s_current_state_reg_38__QN) );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF ( .D(StateRegInput[38]), .CK(
        clk), .Q(Ciphertext[38]), .QN() );
  INV_X1 StateReg_s_current_state_reg_37__U1 ( .A(Ciphertext[37]), .ZN(
        StateReg_s_current_state_reg_37__QN) );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF ( .D(StateRegInput[37]), .CK(
        clk), .Q(Ciphertext[37]), .QN() );
  INV_X1 StateReg_s_current_state_reg_36__U1 ( .A(Ciphertext[36]), .ZN(
        StateReg_s_current_state_reg_36__QN) );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF ( .D(StateRegInput[36]), .CK(
        clk), .Q(Ciphertext[36]), .QN() );
  INV_X1 StateReg_s_current_state_reg_35__U1 ( .A(Ciphertext[35]), .ZN(
        StateReg_s_current_state_reg_35__QN) );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF ( .D(StateRegInput[35]), .CK(
        clk), .Q(Ciphertext[35]), .QN() );
  INV_X1 StateReg_s_current_state_reg_34__U1 ( .A(Ciphertext[34]), .ZN(
        StateReg_s_current_state_reg_34__QN) );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF ( .D(StateRegInput[34]), .CK(
        clk), .Q(Ciphertext[34]), .QN() );
  INV_X1 StateReg_s_current_state_reg_33__U1 ( .A(Ciphertext[33]), .ZN(
        StateReg_s_current_state_reg_33__QN) );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF ( .D(StateRegInput[33]), .CK(
        clk), .Q(Ciphertext[33]), .QN() );
  INV_X1 StateReg_s_current_state_reg_32__U1 ( .A(Ciphertext[32]), .ZN(
        StateReg_s_current_state_reg_32__QN) );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF ( .D(StateRegInput[32]), .CK(
        clk), .Q(Ciphertext[32]), .QN() );
  INV_X1 StateReg_s_current_state_reg_31__U1 ( .A(Ciphertext[31]), .ZN(
        StateReg_s_current_state_reg_31__QN) );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF ( .D(StateRegInput[31]), .CK(
        clk), .Q(Ciphertext[31]), .QN() );
  INV_X1 StateReg_s_current_state_reg_30__U1 ( .A(Ciphertext[30]), .ZN(
        StateReg_s_current_state_reg_30__QN) );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF ( .D(StateRegInput[30]), .CK(
        clk), .Q(Ciphertext[30]), .QN() );
  INV_X1 StateReg_s_current_state_reg_29__U1 ( .A(Ciphertext[29]), .ZN(
        StateReg_s_current_state_reg_29__QN) );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF ( .D(StateRegInput[29]), .CK(
        clk), .Q(Ciphertext[29]), .QN() );
  INV_X1 StateReg_s_current_state_reg_28__U1 ( .A(Ciphertext[28]), .ZN(
        StateReg_s_current_state_reg_28__QN) );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF ( .D(StateRegInput[28]), .CK(
        clk), .Q(Ciphertext[28]), .QN() );
  INV_X1 StateReg_s_current_state_reg_27__U1 ( .A(Ciphertext[27]), .ZN(
        StateReg_s_current_state_reg_27__QN) );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF ( .D(StateRegInput[27]), .CK(
        clk), .Q(Ciphertext[27]), .QN() );
  INV_X1 StateReg_s_current_state_reg_26__U1 ( .A(Ciphertext[26]), .ZN(
        StateReg_s_current_state_reg_26__QN) );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF ( .D(StateRegInput[26]), .CK(
        clk), .Q(Ciphertext[26]), .QN() );
  INV_X1 StateReg_s_current_state_reg_25__U1 ( .A(Ciphertext[25]), .ZN(
        StateReg_s_current_state_reg_25__QN) );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF ( .D(StateRegInput[25]), .CK(
        clk), .Q(Ciphertext[25]), .QN() );
  INV_X1 StateReg_s_current_state_reg_24__U1 ( .A(Ciphertext[24]), .ZN(
        StateReg_s_current_state_reg_24__QN) );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF ( .D(StateRegInput[24]), .CK(
        clk), .Q(Ciphertext[24]), .QN() );
  INV_X1 StateReg_s_current_state_reg_23__U1 ( .A(Ciphertext[23]), .ZN(
        StateReg_s_current_state_reg_23__QN) );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF ( .D(StateRegInput[23]), .CK(
        clk), .Q(Ciphertext[23]), .QN() );
  INV_X1 StateReg_s_current_state_reg_22__U1 ( .A(Ciphertext[22]), .ZN(
        StateReg_s_current_state_reg_22__QN) );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF ( .D(StateRegInput[22]), .CK(
        clk), .Q(Ciphertext[22]), .QN() );
  INV_X1 StateReg_s_current_state_reg_21__U1 ( .A(Ciphertext[21]), .ZN(
        StateReg_s_current_state_reg_21__QN) );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF ( .D(StateRegInput[21]), .CK(
        clk), .Q(Ciphertext[21]), .QN() );
  INV_X1 StateReg_s_current_state_reg_20__U1 ( .A(Ciphertext[20]), .ZN(
        StateReg_s_current_state_reg_20__QN) );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF ( .D(StateRegInput[20]), .CK(
        clk), .Q(Ciphertext[20]), .QN() );
  INV_X1 StateReg_s_current_state_reg_19__U1 ( .A(Ciphertext[19]), .ZN(
        StateReg_s_current_state_reg_19__QN) );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF ( .D(StateRegInput[19]), .CK(
        clk), .Q(Ciphertext[19]), .QN() );
  INV_X1 StateReg_s_current_state_reg_18__U1 ( .A(Ciphertext[18]), .ZN(
        StateReg_s_current_state_reg_18__QN) );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF ( .D(StateRegInput[18]), .CK(
        clk), .Q(Ciphertext[18]), .QN() );
  INV_X1 StateReg_s_current_state_reg_17__U1 ( .A(Ciphertext[17]), .ZN(
        StateReg_s_current_state_reg_17__QN) );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF ( .D(StateRegInput[17]), .CK(
        clk), .Q(Ciphertext[17]), .QN() );
  INV_X1 StateReg_s_current_state_reg_16__U1 ( .A(Ciphertext[16]), .ZN(
        StateReg_s_current_state_reg_16__QN) );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF ( .D(StateRegInput[16]), .CK(
        clk), .Q(Ciphertext[16]), .QN() );
  INV_X1 StateReg_s_current_state_reg_15__U1 ( .A(Ciphertext[15]), .ZN(
        StateReg_s_current_state_reg_15__QN) );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF ( .D(StateRegInput[15]), .CK(
        clk), .Q(Ciphertext[15]), .QN() );
  INV_X1 StateReg_s_current_state_reg_14__U1 ( .A(Ciphertext[14]), .ZN(
        StateReg_s_current_state_reg_14__QN) );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF ( .D(StateRegInput[14]), .CK(
        clk), .Q(Ciphertext[14]), .QN() );
  INV_X1 StateReg_s_current_state_reg_13__U1 ( .A(Ciphertext[13]), .ZN(
        StateReg_s_current_state_reg_13__QN) );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF ( .D(StateRegInput[13]), .CK(
        clk), .Q(Ciphertext[13]), .QN() );
  INV_X1 StateReg_s_current_state_reg_12__U1 ( .A(Ciphertext[12]), .ZN(
        StateReg_s_current_state_reg_12__QN) );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF ( .D(StateRegInput[12]), .CK(
        clk), .Q(Ciphertext[12]), .QN() );
  INV_X1 StateReg_s_current_state_reg_11__U1 ( .A(Ciphertext[11]), .ZN(
        StateReg_s_current_state_reg_11__QN) );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF ( .D(StateRegInput[11]), .CK(
        clk), .Q(Ciphertext[11]), .QN() );
  INV_X1 StateReg_s_current_state_reg_10__U1 ( .A(Ciphertext[10]), .ZN(
        StateReg_s_current_state_reg_10__QN) );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF ( .D(StateRegInput[10]), .CK(
        clk), .Q(Ciphertext[10]), .QN() );
  INV_X1 StateReg_s_current_state_reg_9__U1 ( .A(Ciphertext[9]), .ZN(
        StateReg_s_current_state_reg_9__QN) );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF ( .D(StateRegInput[9]), .CK(clk), .Q(Ciphertext[9]), .QN() );
  INV_X1 StateReg_s_current_state_reg_8__U1 ( .A(Ciphertext[8]), .ZN(
        StateReg_s_current_state_reg_8__QN) );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF ( .D(StateRegInput[8]), .CK(clk), .Q(Ciphertext[8]), .QN() );
  INV_X1 StateReg_s_current_state_reg_7__U1 ( .A(Ciphertext[7]), .ZN(
        StateReg_s_current_state_reg_7__QN) );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF ( .D(StateRegInput[7]), .CK(clk), .Q(Ciphertext[7]), .QN() );
  INV_X1 StateReg_s_current_state_reg_6__U1 ( .A(Ciphertext[6]), .ZN(
        StateReg_s_current_state_reg_6__QN) );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF ( .D(StateRegInput[6]), .CK(clk), .Q(Ciphertext[6]), .QN() );
  INV_X1 StateReg_s_current_state_reg_5__U1 ( .A(Ciphertext[5]), .ZN(
        StateReg_s_current_state_reg_5__QN) );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF ( .D(StateRegInput[5]), .CK(clk), .Q(Ciphertext[5]), .QN() );
  INV_X1 StateReg_s_current_state_reg_4__U1 ( .A(Ciphertext[4]), .ZN(
        StateReg_s_current_state_reg_4__QN) );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF ( .D(StateRegInput[4]), .CK(clk), .Q(Ciphertext[4]), .QN() );
  INV_X1 StateReg_s_current_state_reg_3__U1 ( .A(Ciphertext[3]), .ZN(
        StateReg_s_current_state_reg_3__QN) );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF ( .D(StateRegInput[3]), .CK(clk), .Q(Ciphertext[3]), .QN() );
  INV_X1 StateReg_s_current_state_reg_2__U1 ( .A(Ciphertext[2]), .ZN(
        StateReg_s_current_state_reg_2__QN) );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF ( .D(StateRegInput[2]), .CK(clk), .Q(Ciphertext[2]), .QN() );
  INV_X1 StateReg_s_current_state_reg_1__U1 ( .A(Ciphertext[1]), .ZN(
        StateReg_s_current_state_reg_1__QN) );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF ( .D(StateRegInput[1]), .CK(clk), .Q(Ciphertext[1]), .QN() );
  INV_X1 StateReg_s_current_state_reg_0__U1 ( .A(Ciphertext[0]), .ZN(
        StateReg_s_current_state_reg_0__QN) );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF ( .D(StateRegInput[0]), .CK(clk), .Q(Ciphertext[0]), .QN() );
  INV_X1 SubCellInst_SboxInst_0_U3 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  INV_X1 SubCellInst_SboxInst_0_U1 ( .A(Ciphertext[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1 ( .A(Ciphertext[2]), .B(
        Ciphertext[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1 ( .A(Ciphertext[0]), .B(
        Ciphertext[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1 ( .A(Ciphertext[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1 ( .A(Ciphertext[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_Q1), .ZN(SubCellInst_SboxInst_0_T0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1 ( .A(SubCellInst_SboxInst_0_Q0), .B(
        SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_Q2) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1 ( .A1(Ciphertext[1]), .A2(
        SubCellInst_SboxInst_0_Q2), .ZN(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1 ( .A(Ciphertext[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_Q4), .ZN(SubCellInst_SboxInst_0_T2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1 ( .A(SubCellInst_SboxInst_0_T1), .B(
        SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1 ( .A(SubCellInst_SboxInst_0_XX_2_), 
        .B(SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1 ( .A(SubCellInst_SboxInst_0_Q1), .B(
        SubCellInst_SboxInst_0_Q6), .ZN(SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1 ( .A(SubCellInst_SboxInst_0_L1), .B(
        SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_Q7) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1 ( .A1(SubCellInst_SboxInst_0_Q6), 
        .A2(SubCellInst_SboxInst_0_Q7), .ZN(SubCellInst_SboxInst_0_T3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1 ( .A(Ciphertext[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1 ( .A(SubCellInst_SboxInst_0_L0), .B(
        SubCellInst_SboxInst_0_L2), .Z(SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1 ( .A(SubCellInst_SboxInst_0_L0), .B(
        SubCellInst_SboxInst_0_T3), .Z(ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1 ( .A(SubCellInst_SboxInst_0_XX_2_), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1 ( .A(SubCellInst_SboxInst_0_L3), .B(
        SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1 ( .A(SubCellInst_SboxInst_0_XX_1_), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), 
        .B(SubCellInst_SboxInst_0_YY_3), .ZN(ShiftRowsOutput[5]) );
  INV_X1 SubCellInst_SboxInst_1_U3 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  INV_X1 SubCellInst_SboxInst_1_U1 ( .A(Ciphertext[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1 ( .A(Ciphertext[6]), .B(
        Ciphertext[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1 ( .A(Ciphertext[4]), .B(
        Ciphertext[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1 ( .A(Ciphertext[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1 ( .A(Ciphertext[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_Q1), .ZN(SubCellInst_SboxInst_1_T0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1 ( .A(SubCellInst_SboxInst_1_Q0), .B(
        SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_Q2) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1 ( .A1(Ciphertext[5]), .A2(
        SubCellInst_SboxInst_1_Q2), .ZN(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1 ( .A(Ciphertext[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_Q4), .ZN(SubCellInst_SboxInst_1_T2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1 ( .A(SubCellInst_SboxInst_1_T1), .B(
        SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1 ( .A(SubCellInst_SboxInst_1_XX_2_), 
        .B(SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1 ( .A(SubCellInst_SboxInst_1_Q1), .B(
        SubCellInst_SboxInst_1_Q6), .ZN(SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1 ( .A(SubCellInst_SboxInst_1_L1), .B(
        SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_Q7) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1 ( .A1(SubCellInst_SboxInst_1_Q6), 
        .A2(SubCellInst_SboxInst_1_Q7), .ZN(SubCellInst_SboxInst_1_T3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1 ( .A(Ciphertext[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1 ( .A(SubCellInst_SboxInst_1_L0), .B(
        SubCellInst_SboxInst_1_L2), .Z(SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1 ( .A(SubCellInst_SboxInst_1_L0), .B(
        SubCellInst_SboxInst_1_T3), .Z(ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1 ( .A(SubCellInst_SboxInst_1_XX_2_), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1 ( .A(SubCellInst_SboxInst_1_L3), .B(
        SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1 ( .A(SubCellInst_SboxInst_1_XX_1_), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), 
        .B(SubCellInst_SboxInst_1_YY_3), .ZN(ShiftRowsOutput[9]) );
  INV_X1 SubCellInst_SboxInst_2_U3 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  INV_X1 SubCellInst_SboxInst_2_U1 ( .A(Ciphertext[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1 ( .A(Ciphertext[10]), .B(
        Ciphertext[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1 ( .A(Ciphertext[8]), .B(
        Ciphertext[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1 ( .A(Ciphertext[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1 ( .A(Ciphertext[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_Q1), .ZN(SubCellInst_SboxInst_2_T0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1 ( .A(SubCellInst_SboxInst_2_Q0), .B(
        SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_Q2) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1 ( .A1(Ciphertext[9]), .A2(
        SubCellInst_SboxInst_2_Q2), .ZN(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1 ( .A(Ciphertext[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_Q4), .ZN(SubCellInst_SboxInst_2_T2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1 ( .A(SubCellInst_SboxInst_2_T1), .B(
        SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1 ( .A(SubCellInst_SboxInst_2_XX_2_), 
        .B(SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1 ( .A(SubCellInst_SboxInst_2_Q1), .B(
        SubCellInst_SboxInst_2_Q6), .ZN(SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1 ( .A(SubCellInst_SboxInst_2_L1), .B(
        SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_Q7) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1 ( .A1(SubCellInst_SboxInst_2_Q6), 
        .A2(SubCellInst_SboxInst_2_Q7), .ZN(SubCellInst_SboxInst_2_T3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1 ( .A(Ciphertext[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1 ( .A(SubCellInst_SboxInst_2_L0), .B(
        SubCellInst_SboxInst_2_L2), .Z(SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1 ( .A(SubCellInst_SboxInst_2_L0), .B(
        SubCellInst_SboxInst_2_T3), .Z(ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1 ( .A(SubCellInst_SboxInst_2_XX_2_), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1 ( .A(SubCellInst_SboxInst_2_L3), .B(
        SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1 ( .A(SubCellInst_SboxInst_2_XX_1_), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), 
        .B(SubCellInst_SboxInst_2_YY_3), .ZN(ShiftRowsOutput[13]) );
  INV_X1 SubCellInst_SboxInst_3_U3 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  INV_X1 SubCellInst_SboxInst_3_U1 ( .A(Ciphertext[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1 ( .A(Ciphertext[14]), .B(
        Ciphertext[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1 ( .A(Ciphertext[12]), .B(
        Ciphertext[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1 ( .A(Ciphertext[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1 ( .A(Ciphertext[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_Q1), .ZN(SubCellInst_SboxInst_3_T0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1 ( .A(SubCellInst_SboxInst_3_Q0), .B(
        SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_Q2) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1 ( .A1(Ciphertext[13]), .A2(
        SubCellInst_SboxInst_3_Q2), .ZN(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1 ( .A(Ciphertext[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_Q4), .ZN(SubCellInst_SboxInst_3_T2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1 ( .A(SubCellInst_SboxInst_3_T1), .B(
        SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1 ( .A(SubCellInst_SboxInst_3_XX_2_), 
        .B(SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1 ( .A(SubCellInst_SboxInst_3_Q1), .B(
        SubCellInst_SboxInst_3_Q6), .ZN(SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1 ( .A(SubCellInst_SboxInst_3_L1), .B(
        SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_Q7) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1 ( .A1(SubCellInst_SboxInst_3_Q6), 
        .A2(SubCellInst_SboxInst_3_Q7), .ZN(SubCellInst_SboxInst_3_T3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1 ( .A(Ciphertext[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1 ( .A(SubCellInst_SboxInst_3_L0), .B(
        SubCellInst_SboxInst_3_L2), .Z(SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1 ( .A(SubCellInst_SboxInst_3_L0), .B(
        SubCellInst_SboxInst_3_T3), .Z(ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1 ( .A(SubCellInst_SboxInst_3_XX_2_), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1 ( .A(SubCellInst_SboxInst_3_L3), .B(
        SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1 ( .A(SubCellInst_SboxInst_3_XX_1_), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), 
        .B(SubCellInst_SboxInst_3_YY_3), .ZN(ShiftRowsOutput[1]) );
  INV_X1 SubCellInst_SboxInst_4_U3 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  INV_X1 SubCellInst_SboxInst_4_U1 ( .A(Ciphertext[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1 ( .A(Ciphertext[18]), .B(
        Ciphertext[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1 ( .A(Ciphertext[16]), .B(
        Ciphertext[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1 ( .A(Ciphertext[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1 ( .A(Ciphertext[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_Q1), .ZN(SubCellInst_SboxInst_4_T0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1 ( .A(SubCellInst_SboxInst_4_Q0), .B(
        SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_Q2) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1 ( .A1(Ciphertext[17]), .A2(
        SubCellInst_SboxInst_4_Q2), .ZN(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1 ( .A(Ciphertext[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_Q4), .ZN(SubCellInst_SboxInst_4_T2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1 ( .A(SubCellInst_SboxInst_4_T1), .B(
        SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1 ( .A(SubCellInst_SboxInst_4_XX_2_), 
        .B(SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1 ( .A(SubCellInst_SboxInst_4_Q1), .B(
        SubCellInst_SboxInst_4_Q6), .ZN(SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1 ( .A(SubCellInst_SboxInst_4_L1), .B(
        SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_Q7) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1 ( .A1(SubCellInst_SboxInst_4_Q6), 
        .A2(SubCellInst_SboxInst_4_Q7), .ZN(SubCellInst_SboxInst_4_T3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1 ( .A(Ciphertext[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1 ( .A(SubCellInst_SboxInst_4_L0), .B(
        SubCellInst_SboxInst_4_L2), .Z(SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1 ( .A(SubCellInst_SboxInst_4_L0), .B(
        SubCellInst_SboxInst_4_T3), .Z(ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1 ( .A(SubCellInst_SboxInst_4_XX_2_), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1 ( .A(SubCellInst_SboxInst_4_L3), .B(
        SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1 ( .A(SubCellInst_SboxInst_4_XX_1_), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), 
        .B(SubCellInst_SboxInst_4_YY_3), .ZN(ShiftRowsOutput[25]) );
  INV_X1 SubCellInst_SboxInst_5_U3 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  INV_X1 SubCellInst_SboxInst_5_U1 ( .A(Ciphertext[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1 ( .A(Ciphertext[22]), .B(
        Ciphertext[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1 ( .A(Ciphertext[20]), .B(
        Ciphertext[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1 ( .A(Ciphertext[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1 ( .A(Ciphertext[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_Q1), .ZN(SubCellInst_SboxInst_5_T0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1 ( .A(SubCellInst_SboxInst_5_Q0), .B(
        SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_Q2) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1 ( .A1(Ciphertext[21]), .A2(
        SubCellInst_SboxInst_5_Q2), .ZN(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1 ( .A(Ciphertext[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_Q4), .ZN(SubCellInst_SboxInst_5_T2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1 ( .A(SubCellInst_SboxInst_5_T1), .B(
        SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1 ( .A(SubCellInst_SboxInst_5_XX_2_), 
        .B(SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1 ( .A(SubCellInst_SboxInst_5_Q1), .B(
        SubCellInst_SboxInst_5_Q6), .ZN(SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1 ( .A(SubCellInst_SboxInst_5_L1), .B(
        SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_Q7) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1 ( .A1(SubCellInst_SboxInst_5_Q6), 
        .A2(SubCellInst_SboxInst_5_Q7), .ZN(SubCellInst_SboxInst_5_T3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1 ( .A(Ciphertext[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1 ( .A(SubCellInst_SboxInst_5_L0), .B(
        SubCellInst_SboxInst_5_L2), .Z(SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1 ( .A(SubCellInst_SboxInst_5_L0), .B(
        SubCellInst_SboxInst_5_T3), .Z(ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1 ( .A(SubCellInst_SboxInst_5_XX_2_), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1 ( .A(SubCellInst_SboxInst_5_L3), .B(
        SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1 ( .A(SubCellInst_SboxInst_5_XX_1_), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), 
        .B(SubCellInst_SboxInst_5_YY_3), .ZN(ShiftRowsOutput[29]) );
  INV_X1 SubCellInst_SboxInst_6_U3 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  INV_X1 SubCellInst_SboxInst_6_U1 ( .A(Ciphertext[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1 ( .A(Ciphertext[26]), .B(
        Ciphertext[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1 ( .A(Ciphertext[24]), .B(
        Ciphertext[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1 ( .A(Ciphertext[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1 ( .A(Ciphertext[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_Q1), .ZN(SubCellInst_SboxInst_6_T0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1 ( .A(SubCellInst_SboxInst_6_Q0), .B(
        SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_Q2) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1 ( .A1(Ciphertext[25]), .A2(
        SubCellInst_SboxInst_6_Q2), .ZN(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1 ( .A(Ciphertext[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_Q4), .ZN(SubCellInst_SboxInst_6_T2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1 ( .A(SubCellInst_SboxInst_6_T1), .B(
        SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1 ( .A(SubCellInst_SboxInst_6_XX_2_), 
        .B(SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1 ( .A(SubCellInst_SboxInst_6_Q1), .B(
        SubCellInst_SboxInst_6_Q6), .ZN(SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1 ( .A(SubCellInst_SboxInst_6_L1), .B(
        SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_Q7) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1 ( .A1(SubCellInst_SboxInst_6_Q6), 
        .A2(SubCellInst_SboxInst_6_Q7), .ZN(SubCellInst_SboxInst_6_T3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1 ( .A(Ciphertext[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1 ( .A(SubCellInst_SboxInst_6_L0), .B(
        SubCellInst_SboxInst_6_L2), .Z(SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1 ( .A(SubCellInst_SboxInst_6_L0), .B(
        SubCellInst_SboxInst_6_T3), .Z(ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1 ( .A(SubCellInst_SboxInst_6_XX_2_), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1 ( .A(SubCellInst_SboxInst_6_L3), .B(
        SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1 ( .A(SubCellInst_SboxInst_6_XX_1_), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), 
        .B(SubCellInst_SboxInst_6_YY_3), .ZN(ShiftRowsOutput[17]) );
  INV_X1 SubCellInst_SboxInst_7_U3 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  INV_X1 SubCellInst_SboxInst_7_U1 ( .A(Ciphertext[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1 ( .A(Ciphertext[30]), .B(
        Ciphertext[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1 ( .A(Ciphertext[28]), .B(
        Ciphertext[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1 ( .A(Ciphertext[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1 ( .A(Ciphertext[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_Q1), .ZN(SubCellInst_SboxInst_7_T0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1 ( .A(SubCellInst_SboxInst_7_Q0), .B(
        SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_Q2) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1 ( .A1(Ciphertext[29]), .A2(
        SubCellInst_SboxInst_7_Q2), .ZN(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1 ( .A(Ciphertext[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_Q4), .ZN(SubCellInst_SboxInst_7_T2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1 ( .A(SubCellInst_SboxInst_7_T1), .B(
        SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1 ( .A(SubCellInst_SboxInst_7_XX_2_), 
        .B(SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1 ( .A(SubCellInst_SboxInst_7_Q1), .B(
        SubCellInst_SboxInst_7_Q6), .ZN(SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1 ( .A(SubCellInst_SboxInst_7_L1), .B(
        SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_Q7) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1 ( .A1(SubCellInst_SboxInst_7_Q6), 
        .A2(SubCellInst_SboxInst_7_Q7), .ZN(SubCellInst_SboxInst_7_T3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1 ( .A(Ciphertext[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1 ( .A(SubCellInst_SboxInst_7_L0), .B(
        SubCellInst_SboxInst_7_L2), .Z(SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1 ( .A(SubCellInst_SboxInst_7_L0), .B(
        SubCellInst_SboxInst_7_T3), .Z(ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1 ( .A(SubCellInst_SboxInst_7_XX_2_), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1 ( .A(SubCellInst_SboxInst_7_L3), .B(
        SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1 ( .A(SubCellInst_SboxInst_7_XX_1_), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), 
        .B(SubCellInst_SboxInst_7_YY_3), .ZN(SubCellOutput[29]) );
  INV_X1 SubCellInst_SboxInst_8_U3 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  INV_X1 SubCellInst_SboxInst_8_U1 ( .A(Ciphertext[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1 ( .A(Ciphertext[34]), .B(
        Ciphertext[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1 ( .A(Ciphertext[32]), .B(
        Ciphertext[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1 ( .A(Ciphertext[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1 ( .A(Ciphertext[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_Q1), .ZN(SubCellInst_SboxInst_8_T0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1 ( .A(SubCellInst_SboxInst_8_Q0), .B(
        SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_Q2) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1 ( .A1(Ciphertext[33]), .A2(
        SubCellInst_SboxInst_8_Q2), .ZN(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1 ( .A(Ciphertext[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_Q4), .ZN(SubCellInst_SboxInst_8_T2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1 ( .A(SubCellInst_SboxInst_8_T1), .B(
        SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1 ( .A(SubCellInst_SboxInst_8_XX_2_), 
        .B(SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1 ( .A(SubCellInst_SboxInst_8_Q1), .B(
        SubCellInst_SboxInst_8_Q6), .ZN(SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1 ( .A(SubCellInst_SboxInst_8_L1), .B(
        SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_Q7) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1 ( .A1(SubCellInst_SboxInst_8_Q6), 
        .A2(SubCellInst_SboxInst_8_Q7), .ZN(SubCellInst_SboxInst_8_T3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1 ( .A(Ciphertext[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1 ( .A(SubCellInst_SboxInst_8_L0), .B(
        SubCellInst_SboxInst_8_L2), .Z(SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1 ( .A(SubCellInst_SboxInst_8_L0), .B(
        SubCellInst_SboxInst_8_T3), .Z(AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1 ( .A(SubCellInst_SboxInst_8_XX_2_), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1 ( .A(SubCellInst_SboxInst_8_L3), .B(
        SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1 ( .A(SubCellInst_SboxInst_8_XX_1_), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), 
        .B(SubCellInst_SboxInst_8_YY_3), .ZN(AddRoundConstantOutput[33]) );
  INV_X1 SubCellInst_SboxInst_9_U3 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  INV_X1 SubCellInst_SboxInst_9_U1 ( .A(Ciphertext[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1 ( .A(Ciphertext[38]), .B(
        Ciphertext[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1 ( .A(Ciphertext[36]), .B(
        Ciphertext[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1 ( .A(Ciphertext[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1 ( .A(Ciphertext[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_Q1), .ZN(SubCellInst_SboxInst_9_T0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1 ( .A(SubCellInst_SboxInst_9_Q0), .B(
        SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_Q2) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1 ( .A1(Ciphertext[37]), .A2(
        SubCellInst_SboxInst_9_Q2), .ZN(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1 ( .A(Ciphertext[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_Q4), .ZN(SubCellInst_SboxInst_9_T2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1 ( .A(SubCellInst_SboxInst_9_T1), .B(
        SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1 ( .A(SubCellInst_SboxInst_9_XX_2_), 
        .B(SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1 ( .A(SubCellInst_SboxInst_9_Q1), .B(
        SubCellInst_SboxInst_9_Q6), .ZN(SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1 ( .A(SubCellInst_SboxInst_9_L1), .B(
        SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_Q7) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1 ( .A1(SubCellInst_SboxInst_9_Q6), 
        .A2(SubCellInst_SboxInst_9_Q7), .ZN(SubCellInst_SboxInst_9_T3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1 ( .A(Ciphertext[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1 ( .A(SubCellInst_SboxInst_9_L0), .B(
        SubCellInst_SboxInst_9_L2), .Z(SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1 ( .A(SubCellInst_SboxInst_9_L0), .B(
        SubCellInst_SboxInst_9_T3), .Z(AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1 ( .A(SubCellInst_SboxInst_9_XX_2_), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1 ( .A(SubCellInst_SboxInst_9_L3), .B(
        SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1 ( .A(SubCellInst_SboxInst_9_XX_1_), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), 
        .B(SubCellInst_SboxInst_9_YY_3), .ZN(AddRoundConstantOutput[37]) );
  INV_X1 SubCellInst_SboxInst_10_U3 ( .A(SubCellInst_SboxInst_10_YY_1_), .ZN(
        AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2 ( .A(SubCellInst_SboxInst_10_YY_0_), .ZN(
        AddRoundConstantOutput[42]) );
  INV_X1 SubCellInst_SboxInst_10_U1 ( .A(Ciphertext[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1 ( .A(Ciphertext[42]), .B(
        Ciphertext[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1 ( .A(Ciphertext[40]), .B(
        Ciphertext[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1 ( .A(Ciphertext[41]), .B(
        SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1 ( .A(Ciphertext[41]), .B(
        SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_Q1), .ZN(SubCellInst_SboxInst_10_T0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1 ( .A(SubCellInst_SboxInst_10_Q0), 
        .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_Q2) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1 ( .A1(Ciphertext[41]), .A2(
        SubCellInst_SboxInst_10_Q2), .ZN(SubCellInst_SboxInst_10_T1) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1 ( .A(Ciphertext[41]), .B(
        SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_Q4), .ZN(SubCellInst_SboxInst_10_T2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1 ( .A(SubCellInst_SboxInst_10_T1), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1 ( .A(SubCellInst_SboxInst_10_XX_2_), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1 ( .A(SubCellInst_SboxInst_10_Q1), 
        .B(SubCellInst_SboxInst_10_Q6), .ZN(SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1 ( .A(SubCellInst_SboxInst_10_L1), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_Q7) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1 ( .A1(SubCellInst_SboxInst_10_Q6), 
        .A2(SubCellInst_SboxInst_10_Q7), .ZN(SubCellInst_SboxInst_10_T3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1 ( .A(Ciphertext[41]), .B(
        SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1 ( .A(SubCellInst_SboxInst_10_L0), 
        .B(SubCellInst_SboxInst_10_L2), .Z(SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1 ( .A(SubCellInst_SboxInst_10_L0), 
        .B(SubCellInst_SboxInst_10_T3), .Z(AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1 ( .A(SubCellInst_SboxInst_10_XX_2_), 
        .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1 ( .A(SubCellInst_SboxInst_10_L3), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1 ( .A(SubCellInst_SboxInst_10_XX_1_), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_10_YY_1_), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  INV_X1 SubCellInst_SboxInst_11_U3 ( .A(SubCellInst_SboxInst_11_YY_1_), .ZN(
        SubCellOutput[47]) );
  INV_X1 SubCellInst_SboxInst_11_U2 ( .A(SubCellInst_SboxInst_11_YY_0_), .ZN(
        SubCellOutput[46]) );
  INV_X1 SubCellInst_SboxInst_11_U1 ( .A(Ciphertext[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1 ( .A(Ciphertext[46]), .B(
        Ciphertext[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1 ( .A(Ciphertext[44]), .B(
        Ciphertext[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1 ( .A(Ciphertext[45]), .B(
        SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1 ( .A(Ciphertext[45]), .B(
        SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_Q1), .ZN(SubCellInst_SboxInst_11_T0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1 ( .A(SubCellInst_SboxInst_11_Q0), 
        .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_Q2) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1 ( .A1(Ciphertext[45]), .A2(
        SubCellInst_SboxInst_11_Q2), .ZN(SubCellInst_SboxInst_11_T1) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1 ( .A(Ciphertext[45]), .B(
        SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_Q4), .ZN(SubCellInst_SboxInst_11_T2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1 ( .A(SubCellInst_SboxInst_11_T1), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1 ( .A(SubCellInst_SboxInst_11_XX_2_), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1 ( .A(SubCellInst_SboxInst_11_Q1), 
        .B(SubCellInst_SboxInst_11_Q6), .ZN(SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1 ( .A(SubCellInst_SboxInst_11_L1), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_Q7) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1 ( .A1(SubCellInst_SboxInst_11_Q6), 
        .A2(SubCellInst_SboxInst_11_Q7), .ZN(SubCellInst_SboxInst_11_T3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1 ( .A(Ciphertext[45]), .B(
        SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1 ( .A(SubCellInst_SboxInst_11_L0), 
        .B(SubCellInst_SboxInst_11_L2), .Z(SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1 ( .A(SubCellInst_SboxInst_11_L0), 
        .B(SubCellInst_SboxInst_11_T3), .Z(SubCellOutput[44]) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1 ( .A(SubCellInst_SboxInst_11_XX_2_), 
        .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1 ( .A(SubCellInst_SboxInst_11_L3), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1 ( .A(SubCellInst_SboxInst_11_XX_1_), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_11_YY_1_), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput[45]) );
  INV_X1 SubCellInst_SboxInst_12_U3 ( .A(SubCellInst_SboxInst_12_YY_1_), .ZN(
        AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2 ( .A(SubCellInst_SboxInst_12_YY_0_), .ZN(
        AddRoundConstantOutput[50]) );
  INV_X1 SubCellInst_SboxInst_12_U1 ( .A(Ciphertext[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1 ( .A(Ciphertext[50]), .B(
        Ciphertext[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1 ( .A(Ciphertext[48]), .B(
        Ciphertext[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1 ( .A(Ciphertext[49]), .B(
        SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1 ( .A(Ciphertext[49]), .B(
        SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_Q1), .ZN(SubCellInst_SboxInst_12_T0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1 ( .A(SubCellInst_SboxInst_12_Q0), 
        .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_Q2) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1 ( .A1(Ciphertext[49]), .A2(
        SubCellInst_SboxInst_12_Q2), .ZN(SubCellInst_SboxInst_12_T1) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1 ( .A(Ciphertext[49]), .B(
        SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_Q4), .ZN(SubCellInst_SboxInst_12_T2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1 ( .A(SubCellInst_SboxInst_12_T1), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1 ( .A(SubCellInst_SboxInst_12_XX_2_), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1 ( .A(SubCellInst_SboxInst_12_Q1), 
        .B(SubCellInst_SboxInst_12_Q6), .ZN(SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1 ( .A(SubCellInst_SboxInst_12_L1), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_Q7) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1 ( .A1(SubCellInst_SboxInst_12_Q6), 
        .A2(SubCellInst_SboxInst_12_Q7), .ZN(SubCellInst_SboxInst_12_T3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1 ( .A(Ciphertext[49]), .B(
        SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1 ( .A(SubCellInst_SboxInst_12_L0), 
        .B(SubCellInst_SboxInst_12_L2), .Z(SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1 ( .A(SubCellInst_SboxInst_12_L0), 
        .B(SubCellInst_SboxInst_12_T3), .Z(AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1 ( .A(SubCellInst_SboxInst_12_XX_2_), 
        .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1 ( .A(SubCellInst_SboxInst_12_L3), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1 ( .A(SubCellInst_SboxInst_12_XX_1_), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_12_YY_1_), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  INV_X1 SubCellInst_SboxInst_13_U3 ( .A(SubCellInst_SboxInst_13_YY_1_), .ZN(
        AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2 ( .A(SubCellInst_SboxInst_13_YY_0_), .ZN(
        AddRoundConstantOutput[54]) );
  INV_X1 SubCellInst_SboxInst_13_U1 ( .A(Ciphertext[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1 ( .A(Ciphertext[54]), .B(
        Ciphertext[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1 ( .A(Ciphertext[52]), .B(
        Ciphertext[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1 ( .A(Ciphertext[53]), .B(
        SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1 ( .A(Ciphertext[53]), .B(
        SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_Q1), .ZN(SubCellInst_SboxInst_13_T0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1 ( .A(SubCellInst_SboxInst_13_Q0), 
        .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_Q2) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1 ( .A1(Ciphertext[53]), .A2(
        SubCellInst_SboxInst_13_Q2), .ZN(SubCellInst_SboxInst_13_T1) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1 ( .A(Ciphertext[53]), .B(
        SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_Q4), .ZN(SubCellInst_SboxInst_13_T2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1 ( .A(SubCellInst_SboxInst_13_T1), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1 ( .A(SubCellInst_SboxInst_13_XX_2_), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1 ( .A(SubCellInst_SboxInst_13_Q1), 
        .B(SubCellInst_SboxInst_13_Q6), .ZN(SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1 ( .A(SubCellInst_SboxInst_13_L1), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_Q7) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1 ( .A1(SubCellInst_SboxInst_13_Q6), 
        .A2(SubCellInst_SboxInst_13_Q7), .ZN(SubCellInst_SboxInst_13_T3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1 ( .A(Ciphertext[53]), .B(
        SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1 ( .A(SubCellInst_SboxInst_13_L0), 
        .B(SubCellInst_SboxInst_13_L2), .Z(SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1 ( .A(SubCellInst_SboxInst_13_L0), 
        .B(SubCellInst_SboxInst_13_T3), .Z(AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1 ( .A(SubCellInst_SboxInst_13_XX_2_), 
        .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1 ( .A(SubCellInst_SboxInst_13_L3), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1 ( .A(SubCellInst_SboxInst_13_XX_1_), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_13_YY_1_), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  INV_X1 SubCellInst_SboxInst_14_U3 ( .A(SubCellInst_SboxInst_14_YY_1_), .ZN(
        AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2 ( .A(SubCellInst_SboxInst_14_YY_0_), .ZN(
        AddRoundConstantOutput[58]) );
  INV_X1 SubCellInst_SboxInst_14_U1 ( .A(Ciphertext[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1 ( .A(Ciphertext[58]), .B(
        Ciphertext[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1 ( .A(Ciphertext[56]), .B(
        Ciphertext[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1 ( .A(Ciphertext[57]), .B(
        SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1 ( .A(Ciphertext[57]), .B(
        SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_Q1), .ZN(SubCellInst_SboxInst_14_T0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1 ( .A(SubCellInst_SboxInst_14_Q0), 
        .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_Q2) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1 ( .A1(Ciphertext[57]), .A2(
        SubCellInst_SboxInst_14_Q2), .ZN(SubCellInst_SboxInst_14_T1) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1 ( .A(Ciphertext[57]), .B(
        SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_Q4), .ZN(SubCellInst_SboxInst_14_T2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1 ( .A(SubCellInst_SboxInst_14_T1), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1 ( .A(SubCellInst_SboxInst_14_XX_2_), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1 ( .A(SubCellInst_SboxInst_14_Q1), 
        .B(SubCellInst_SboxInst_14_Q6), .ZN(SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1 ( .A(SubCellInst_SboxInst_14_L1), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_Q7) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1 ( .A1(SubCellInst_SboxInst_14_Q6), 
        .A2(SubCellInst_SboxInst_14_Q7), .ZN(SubCellInst_SboxInst_14_T3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1 ( .A(Ciphertext[57]), .B(
        SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1 ( .A(SubCellInst_SboxInst_14_L0), 
        .B(SubCellInst_SboxInst_14_L2), .Z(SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1 ( .A(SubCellInst_SboxInst_14_L0), 
        .B(SubCellInst_SboxInst_14_T3), .Z(AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1 ( .A(SubCellInst_SboxInst_14_XX_2_), 
        .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1 ( .A(SubCellInst_SboxInst_14_L3), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1 ( .A(SubCellInst_SboxInst_14_XX_1_), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_14_YY_1_), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  INV_X1 SubCellInst_SboxInst_15_U3 ( .A(SubCellInst_SboxInst_15_YY_1_), .ZN(
        SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2 ( .A(SubCellInst_SboxInst_15_YY_0_), .ZN(
        SubCellOutput[62]) );
  INV_X1 SubCellInst_SboxInst_15_U1 ( .A(Ciphertext[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1 ( .A(Ciphertext[62]), .B(
        Ciphertext[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1 ( .A(Ciphertext[60]), .B(
        Ciphertext[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1 ( .A(Ciphertext[61]), .B(
        SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1 ( .A(Ciphertext[61]), .B(
        SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_Q1), .ZN(SubCellInst_SboxInst_15_T0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1 ( .A(SubCellInst_SboxInst_15_Q0), 
        .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_Q2) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1 ( .A1(Ciphertext[61]), .A2(
        SubCellInst_SboxInst_15_Q2), .ZN(SubCellInst_SboxInst_15_T1) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1 ( .A(Ciphertext[61]), .B(
        SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_Q4), .ZN(SubCellInst_SboxInst_15_T2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1 ( .A(SubCellInst_SboxInst_15_T1), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1 ( .A(SubCellInst_SboxInst_15_XX_2_), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_Q6) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1 ( .A(SubCellInst_SboxInst_15_Q1), 
        .B(SubCellInst_SboxInst_15_Q6), .ZN(SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1 ( .A(SubCellInst_SboxInst_15_L1), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_Q7) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1 ( .A1(SubCellInst_SboxInst_15_Q6), 
        .A2(SubCellInst_SboxInst_15_Q7), .ZN(SubCellInst_SboxInst_15_T3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1 ( .A(Ciphertext[61]), .B(
        SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1 ( .A(SubCellInst_SboxInst_15_L0), 
        .B(SubCellInst_SboxInst_15_L2), .Z(SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1 ( .A(SubCellInst_SboxInst_15_L0), 
        .B(SubCellInst_SboxInst_15_T3), .Z(SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1 ( .A(SubCellInst_SboxInst_15_XX_2_), 
        .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1 ( .A(SubCellInst_SboxInst_15_L3), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1 ( .A(SubCellInst_SboxInst_15_XX_1_), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_YY_0_) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1 ( .A(
        SubCellInst_SboxInst_15_YY_1_), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  INV_X1 AddConstXOR_U2 ( .A(SubCellOutput[29]), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(FSMUpdate[1]), .ZN(
        AddRoundConstantOutput[60]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(FSM[1]), .ZN(
        AddRoundConstantOutput[61]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(FSMUpdate[3]), .ZN(
        AddRoundConstantOutput[62]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(FSMUpdate[4]), .ZN(
        AddRoundConstantOutput[63]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(FSM[4]), .ZN(
        AddRoundConstantOutput[44]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .A(1'b0), .B(
        SubCellOutput[44]), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(FSM[5]), .ZN(
        AddRoundConstantOutput[45]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .A(1'b0), .B(
        SubCellOutput[45]), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .A(1'b0), .B(
        SubCellOutput[46]), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .A(1'b0), .B(
        SubCellOutput[47]), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(
        TweakeyGeneration_key_Feedback[0]), .ZN(ShiftRowsOutput[44]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(
        TweakeyGeneration_key_Feedback[1]), .ZN(ShiftRowsOutput[45]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(
        TweakeyGeneration_key_Feedback[2]), .ZN(ShiftRowsOutput[46]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(
        TweakeyGeneration_key_Feedback[3]), .ZN(ShiftRowsOutput[47]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(
        TweakeyGeneration_key_Feedback[4]), .ZN(ShiftRowsOutput[32]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(
        TweakeyGeneration_key_Feedback[5]), .ZN(ShiftRowsOutput[33]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(
        TweakeyGeneration_key_Feedback[6]), .ZN(ShiftRowsOutput[34]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(
        TweakeyGeneration_key_Feedback[7]), .ZN(ShiftRowsOutput[35]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(
        TweakeyGeneration_key_Feedback[8]), .ZN(ShiftRowsOutput[36]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(
        TweakeyGeneration_key_Feedback[9]), .ZN(ShiftRowsOutput[37]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(
        TweakeyGeneration_key_Feedback[10]), .ZN(ShiftRowsOutput[38]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(
        TweakeyGeneration_key_Feedback[11]), .ZN(ShiftRowsOutput[39]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(
        TweakeyGeneration_key_Feedback[12]), .ZN(ShiftRowsOutput[40]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(
        TweakeyGeneration_key_Feedback[13]), .ZN(ShiftRowsOutput[41]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(
        TweakeyGeneration_key_Feedback[14]), .ZN(ShiftRowsOutput[42]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(
        TweakeyGeneration_key_Feedback[15]), .ZN(ShiftRowsOutput[43]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(
        TweakeyGeneration_key_Feedback[16]), .ZN(MCOutput[32]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(
        TweakeyGeneration_key_Feedback[17]), .ZN(MCOutput[33]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(
        TweakeyGeneration_key_Feedback[18]), .ZN(MCOutput[34]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(
        TweakeyGeneration_key_Feedback[19]), .ZN(MCOutput[35]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(
        TweakeyGeneration_key_Feedback[20]), .ZN(MCOutput[36]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(
        TweakeyGeneration_key_Feedback[21]), .ZN(MCOutput[37]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(
        TweakeyGeneration_key_Feedback[22]), .ZN(MCOutput[38]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(
        TweakeyGeneration_key_Feedback[23]), .ZN(MCOutput[39]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(
        TweakeyGeneration_key_Feedback[24]), .ZN(MCOutput[40]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(
        TweakeyGeneration_key_Feedback[25]), .ZN(MCOutput[41]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(
        TweakeyGeneration_key_Feedback[26]), .ZN(MCOutput[42]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(
        TweakeyGeneration_key_Feedback[27]), .ZN(MCOutput[43]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(
        TweakeyGeneration_key_Feedback[28]), .ZN(MCOutput[44]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(
        TweakeyGeneration_key_Feedback[29]), .ZN(MCOutput[45]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(
        TweakeyGeneration_key_Feedback[30]), .ZN(MCOutput[46]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(
        TweakeyGeneration_key_Feedback[31]), .ZN(MCOutput[47]) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3 ( .A(MCInst_MCR0_XORInst_0_0_n2), .B(
        MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[32]), .Z(
        MCInst_MCR0_XORInst_0_0_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3 ( .A(MCInst_MCR0_XORInst_0_1_n2), .B(
        MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[33]), .Z(
        MCInst_MCR0_XORInst_0_1_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3 ( .A(MCInst_MCR0_XORInst_0_2_n2), .B(
        MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[34]), .Z(
        MCInst_MCR0_XORInst_0_2_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3 ( .A(MCInst_MCR0_XORInst_0_3_n2), .B(
        MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[35]), .Z(
        MCInst_MCR0_XORInst_0_3_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3 ( .A(MCInst_MCR0_XORInst_1_0_n2), .B(
        MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[36]), .Z(
        MCInst_MCR0_XORInst_1_0_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3 ( .A(MCInst_MCR0_XORInst_1_1_n2), .B(
        MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[37]), .Z(
        MCInst_MCR0_XORInst_1_1_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3 ( .A(MCInst_MCR0_XORInst_1_2_n2), .B(
        MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[38]), .Z(
        MCInst_MCR0_XORInst_1_2_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3 ( .A(MCInst_MCR0_XORInst_1_3_n2), .B(
        MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[39]), .Z(
        MCInst_MCR0_XORInst_1_3_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3 ( .A(MCInst_MCR0_XORInst_2_0_n2), .B(
        MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[40]), .Z(
        MCInst_MCR0_XORInst_2_0_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3 ( .A(MCInst_MCR0_XORInst_2_1_n2), .B(
        MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[41]), .Z(
        MCInst_MCR0_XORInst_2_1_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3 ( .A(MCInst_MCR0_XORInst_2_2_n2), .B(
        MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[42]), .Z(
        MCInst_MCR0_XORInst_2_2_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3 ( .A(MCInst_MCR0_XORInst_2_3_n2), .B(
        MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[43]), .Z(
        MCInst_MCR0_XORInst_2_3_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3 ( .A(MCInst_MCR0_XORInst_3_0_n2), .B(
        MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[44]), .Z(
        MCInst_MCR0_XORInst_3_0_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3 ( .A(MCInst_MCR0_XORInst_3_1_n2), .B(
        MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[45]), .Z(
        MCInst_MCR0_XORInst_3_1_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3 ( .A(MCInst_MCR0_XORInst_3_2_n2), .B(
        MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[46]), .Z(
        MCInst_MCR0_XORInst_3_2_n2) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3 ( .A(MCInst_MCR0_XORInst_3_3_n2), .B(
        MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[47]), .Z(
        MCInst_MCR0_XORInst_3_3_n2) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2 ( .A(MCInst_MCR2_XORInst_0_0_n1), .B(
        ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1 ( .A(1'b0), .B(ShiftRowsOutput[32]), 
        .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2 ( .A(MCInst_MCR2_XORInst_0_1_n1), .B(
        ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1 ( .A(1'b0), .B(ShiftRowsOutput[33]), 
        .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2 ( .A(MCInst_MCR2_XORInst_0_2_n1), .B(
        ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1 ( .A(1'b0), .B(ShiftRowsOutput[34]), 
        .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2 ( .A(MCInst_MCR2_XORInst_0_3_n1), .B(
        ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1 ( .A(1'b0), .B(ShiftRowsOutput[35]), 
        .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2 ( .A(MCInst_MCR2_XORInst_1_0_n1), .B(
        ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1 ( .A(1'b0), .B(ShiftRowsOutput[36]), 
        .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2 ( .A(MCInst_MCR2_XORInst_1_1_n1), .B(
        ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1 ( .A(1'b0), .B(ShiftRowsOutput[37]), 
        .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2 ( .A(MCInst_MCR2_XORInst_1_2_n1), .B(
        ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1 ( .A(1'b0), .B(ShiftRowsOutput[38]), 
        .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2 ( .A(MCInst_MCR2_XORInst_1_3_n1), .B(
        ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1 ( .A(1'b0), .B(ShiftRowsOutput[39]), 
        .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2 ( .A(MCInst_MCR2_XORInst_2_0_n1), .B(
        ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1 ( .A(1'b0), .B(ShiftRowsOutput[40]), 
        .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2 ( .A(MCInst_MCR2_XORInst_2_1_n1), .B(
        ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1 ( .A(1'b0), .B(ShiftRowsOutput[41]), 
        .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2 ( .A(MCInst_MCR2_XORInst_2_2_n1), .B(
        ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1 ( .A(1'b0), .B(ShiftRowsOutput[42]), 
        .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2 ( .A(MCInst_MCR2_XORInst_2_3_n1), .B(
        ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1 ( .A(1'b0), .B(ShiftRowsOutput[43]), 
        .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2 ( .A(MCInst_MCR2_XORInst_3_0_n1), .B(
        ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1 ( .A(1'b0), .B(ShiftRowsOutput[44]), 
        .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2 ( .A(MCInst_MCR2_XORInst_3_1_n1), .B(
        ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1 ( .A(1'b0), .B(ShiftRowsOutput[45]), 
        .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2 ( .A(MCInst_MCR2_XORInst_3_2_n1), .B(
        ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1 ( .A(1'b0), .B(ShiftRowsOutput[46]), 
        .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2 ( .A(MCInst_MCR2_XORInst_3_3_n1), .B(
        ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1 ( .A(1'b0), .B(ShiftRowsOutput[47]), 
        .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2 ( .A(MCInst_MCR3_XORInst_0_0_n1), .B(
        ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[32]), .ZN(
        MCInst_MCR3_XORInst_0_0_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2 ( .A(MCInst_MCR3_XORInst_0_1_n1), .B(
        ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[33]), .ZN(
        MCInst_MCR3_XORInst_0_1_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2 ( .A(MCInst_MCR3_XORInst_0_2_n1), .B(
        ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[34]), .ZN(
        MCInst_MCR3_XORInst_0_2_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2 ( .A(MCInst_MCR3_XORInst_0_3_n1), .B(
        ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[35]), .ZN(
        MCInst_MCR3_XORInst_0_3_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2 ( .A(MCInst_MCR3_XORInst_1_0_n1), .B(
        ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[36]), .ZN(
        MCInst_MCR3_XORInst_1_0_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2 ( .A(MCInst_MCR3_XORInst_1_1_n1), .B(
        ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[37]), .ZN(
        MCInst_MCR3_XORInst_1_1_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2 ( .A(MCInst_MCR3_XORInst_1_2_n1), .B(
        ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[38]), .ZN(
        MCInst_MCR3_XORInst_1_2_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2 ( .A(MCInst_MCR3_XORInst_1_3_n1), .B(
        ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[39]), .ZN(
        MCInst_MCR3_XORInst_1_3_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2 ( .A(MCInst_MCR3_XORInst_2_0_n1), .B(
        ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[40]), .ZN(
        MCInst_MCR3_XORInst_2_0_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2 ( .A(MCInst_MCR3_XORInst_2_1_n1), .B(
        ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[41]), .ZN(
        MCInst_MCR3_XORInst_2_1_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2 ( .A(MCInst_MCR3_XORInst_2_2_n1), .B(
        ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[42]), .ZN(
        MCInst_MCR3_XORInst_2_2_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2 ( .A(MCInst_MCR3_XORInst_2_3_n1), .B(
        ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[43]), .ZN(
        MCInst_MCR3_XORInst_2_3_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2 ( .A(MCInst_MCR3_XORInst_3_0_n1), .B(
        ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[44]), .ZN(
        MCInst_MCR3_XORInst_3_0_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2 ( .A(MCInst_MCR3_XORInst_3_1_n1), .B(
        ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[45]), .ZN(
        MCInst_MCR3_XORInst_3_1_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2 ( .A(MCInst_MCR3_XORInst_3_2_n1), .B(
        ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[46]), .ZN(
        MCInst_MCR3_XORInst_3_2_n1) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2 ( .A(MCInst_MCR3_XORInst_3_3_n1), .B(
        ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[47]), .ZN(
        MCInst_MCR3_XORInst_3_3_n1) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_63__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[63]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_62__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[62]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_61__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[61]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_60__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[60]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_59__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[59]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_58__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[58]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_57__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[57]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_56__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[56]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_55__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[55]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_54__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[54]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_53__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[53]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_52__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[52]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_51__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[51]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_50__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[50]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_49__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[49]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_48__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[48]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_47__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[47]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_46__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[46]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_45__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[45]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_44__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[44]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_43__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[43]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_42__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[42]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_41__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[41]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_40__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[40]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_39__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[39]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_38__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[38]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_37__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[37]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_36__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[36]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_35__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[35]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_34__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[34]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_33__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[33]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_32__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[32]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_31__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[31]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_30__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[30]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_29__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[29]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_28__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[28]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_27__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[27]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_26__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[26]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_25__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[25]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_24__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[24]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_23__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[23]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_22__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[22]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_21__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[21]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_20__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[20]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_19__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[19]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_18__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[18]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_17__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[17]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_16__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[16]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_15__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[15]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_14__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[14]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_13__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[13]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_12__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[12]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_11__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[11]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_10__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[10]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_9__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[9]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_8__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[8]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_7__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[7]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_6__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[6]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_5__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[5]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_4__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[4]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_3__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[3]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_2__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[2]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_1__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[1]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  INV_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .ZN(
        TweakeyGeneration_StateReg_s_current_state_reg_0__QN) );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .D(
        TweakeyGeneration_StateRegInput[0]), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  MUX2_X1 FSMMUX_MUXInst_0_U1 ( .A(FSMUpdate[0]), .B(1'b1), .S(rst), .Z(
        FSMSelected[0]) );
  MUX2_X1 FSMMUX_MUXInst_1_U1 ( .A(FSMUpdate[1]), .B(1'b0), .S(rst), .Z(
        FSMSelected[1]) );
  MUX2_X1 FSMMUX_MUXInst_2_U1 ( .A(FSMUpdate[2]), .B(1'b0), .S(rst), .Z(
        FSMSelected[2]) );
  MUX2_X1 FSMMUX_MUXInst_3_U1 ( .A(FSMUpdate[3]), .B(1'b0), .S(rst), .Z(
        FSMSelected[3]) );
  MUX2_X1 FSMMUX_MUXInst_4_U1 ( .A(FSMUpdate[4]), .B(1'b0), .S(rst), .Z(
        FSMSelected[4]) );
  MUX2_X1 FSMMUX_MUXInst_5_U1 ( .A(FSMUpdate[5]), .B(1'b0), .S(rst), .Z(
        FSMSelected[5]) );
  INV_X1 FSMReg_s_current_state_reg_5__U1 ( .A(FSM[5]), .ZN(
        FSMReg_s_current_state_reg_5__QN) );
  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(FSMSelected[5]), .CK(clk), 
        .Q(FSM[5]), .QN() );
  INV_X1 FSMReg_s_current_state_reg_4__U1 ( .A(FSM[4]), .ZN(
        FSMReg_s_current_state_reg_4__QN) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(FSMSelected[4]), .CK(clk), 
        .Q(FSM[4]), .QN() );
  INV_X1 FSMReg_s_current_state_reg_3__U1 ( .A(FSMUpdate[4]), .ZN(
        FSMReg_s_current_state_reg_3__QN) );
  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(FSMSelected[3]), .CK(clk), 
        .Q(FSMUpdate[4]), .QN() );
  INV_X1 FSMReg_s_current_state_reg_2__U1 ( .A(FSMUpdate[3]), .ZN(
        FSMReg_s_current_state_reg_2__QN) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(FSMSelected[2]), .CK(clk), 
        .Q(FSMUpdate[3]), .QN() );
  INV_X1 FSMReg_s_current_state_reg_1__U1 ( .A(FSM[1]), .ZN(
        FSMReg_s_current_state_reg_1__QN) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(FSMSelected[1]), .CK(clk), 
        .Q(FSM[1]), .QN() );
  INV_X1 FSMReg_s_current_state_reg_0__U1 ( .A(FSMUpdate[1]), .ZN(
        FSMReg_s_current_state_reg_0__QN) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(FSMSelected[0]), .CK(clk), 
        .Q(FSMUpdate[1]), .QN() );
  MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .A(
        FSMUpdateInst_StateUpdateInst_0_n4), .B(FSM[5]), .S(FSM[4]), .Z(
        FSMUpdate[0]) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1(FSM[5]), .A2(
        FSMUpdateInst_StateUpdateInst_0_n3), .ZN(
        FSMUpdateInst_StateUpdateInst_0_n4) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1(
        FSMUpdateInst_StateUpdateInst_0_n2), .A2(
        FSMUpdateInst_StateUpdateInst_0_n1), .ZN(
        FSMUpdateInst_StateUpdateInst_0_n3) );
  NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1(FSMUpdate[3]), .A2(
        FSMUpdate[4]), .ZN(FSMUpdateInst_StateUpdateInst_0_n1) );
  AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1(FSMUpdate[1]), .A2(FSM[1]), 
        .ZN(FSMUpdateInst_StateUpdateInst_0_n2) );
  AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1(
        FSMUpdateInst_StateUpdateInst_2_n4), .A2(FSM[1]), .ZN(FSMUpdate[2]) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1(
        FSMUpdateInst_StateUpdateInst_2_n3), .A2(FSM[5]), .ZN(
        FSMUpdateInst_StateUpdateInst_2_n4) );
  NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1(FSM[4]), .A2(
        FSMUpdateInst_StateUpdateInst_2_n2), .ZN(
        FSMUpdateInst_StateUpdateInst_2_n3) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1(FSMUpdate[1]), .A2(
        FSMUpdateInst_StateUpdateInst_2_n1), .ZN(
        FSMUpdateInst_StateUpdateInst_2_n2) );
  NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1(FSMUpdate[3]), .A2(
        FSMUpdate[4]), .ZN(FSMUpdateInst_StateUpdateInst_2_n1) );
  OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1(FSM[4]), .A2(
        FSMUpdateInst_StateUpdateInst_5_n4), .ZN(FSMUpdate[5]) );
  NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1(FSMUpdate[4]), .A2(
        FSMUpdateInst_StateUpdateInst_5_n3), .ZN(
        FSMUpdateInst_StateUpdateInst_5_n4) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1(FSM[5]), .A2(
        FSMUpdateInst_StateUpdateInst_5_n2), .ZN(
        FSMUpdateInst_StateUpdateInst_5_n3) );
  NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1(FSMUpdate[3]), .A2(
        FSMUpdateInst_StateUpdateInst_5_n1), .ZN(
        FSMUpdateInst_StateUpdateInst_5_n2) );
  NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1(FSMUpdate[1]), .A2(FSM[1]), 
        .ZN(FSMUpdateInst_StateUpdateInst_5_n1) );
  NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1(FSMSignalsInst_doneInst_n5), .A2(
        FSMSignalsInst_doneInst_n4), .ZN(done) );
  NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1(FSM[4]), .A2(FSM[5]), .ZN(
        FSMSignalsInst_doneInst_n4) );
  NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1(FSMSignalsInst_doneInst_n3), .A2(
        FSMSignalsInst_doneInst_n2), .ZN(FSMSignalsInst_doneInst_n5) );
  NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1(FSMUpdate[4]), .A2(
        FSMSignalsInst_doneInst_n1), .ZN(FSMSignalsInst_doneInst_n2) );
  INV_X1 FSMSignalsInst_doneInst_U2 ( .A(FSMUpdate[1]), .ZN(
        FSMSignalsInst_doneInst_n1) );
  NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1(FSM[1]), .A2(FSMUpdate[3]), .ZN(
        FSMSignalsInst_doneInst_n3) );
endmodule

