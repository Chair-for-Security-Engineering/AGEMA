module LED ( IN_plaintext, IN_key, IN_reset, CLK, OUT_ciphertext, OUT_done );
 (* AGEMA = "secure" *) input [63:0]  IN_plaintext;
 (* AGEMA = "secure" *) input [127:0] IN_key;
 (* AGEMA = "reset" *)  input IN_reset;
 (* AGEMA = "clock" *)  input CLK;
 
  output [63:0] OUT_ciphertext;
  (* AGEMA = "control" *) output OUT_done;

  wire   n15, n14, n16, n17, n18, n19, n20, LED_128_Instance_n34,
         LED_128_Instance_n33, LED_128_Instance_n32, LED_128_Instance_n23,
         LED_128_Instance_n21, LED_128_Instance_n20, LED_128_Instance_n19,
         LED_128_Instance_n18, LED_128_Instance_n17, LED_128_Instance_n16,
         LED_128_Instance_n15, LED_128_Instance_n14, LED_128_Instance_n13,
         LED_128_Instance_n12, LED_128_Instance_n11, LED_128_Instance_n10,
         LED_128_Instance_n2, LED_128_Instance_n1, LED_128_Instance_n27,
         LED_128_Instance_N9, LED_128_Instance_n28, LED_128_Instance_N8,
         LED_128_Instance_n30, LED_128_Instance_N7, LED_128_Instance_n5,
         LED_128_Instance_N6, LED_128_Instance_n29, LED_128_Instance_N5,
         LED_128_Instance_n6, LED_128_Instance_N4, LED_128_Instance_n24,
         LED_128_Instance_N13, LED_128_Instance_n25, LED_128_Instance_N12,
         LED_128_Instance_n8, LED_128_Instance_n26, LED_128_Instance_N11,
         LED_128_Instance_n4, LED_128_Instance_N10, LED_128_Instance_n31,
         LED_128_Instance_addroundkey_out_0_,
         LED_128_Instance_addroundkey_out_1_,
         LED_128_Instance_addroundkey_out_2_,
         LED_128_Instance_addroundkey_out_3_,
         LED_128_Instance_addroundkey_out_4_,
         LED_128_Instance_addroundkey_out_5_,
         LED_128_Instance_addroundkey_out_6_,
         LED_128_Instance_addroundkey_out_16_,
         LED_128_Instance_addroundkey_out_17_,
         LED_128_Instance_addroundkey_out_18_,
         LED_128_Instance_addroundkey_out_19_,
         LED_128_Instance_addroundkey_out_20_,
         LED_128_Instance_addroundkey_out_21_,
         LED_128_Instance_addroundkey_out_22_,
         LED_128_Instance_addroundkey_out_32_,
         LED_128_Instance_addroundkey_out_33_,
         LED_128_Instance_addroundkey_out_34_,
         LED_128_Instance_addroundkey_out_35_,
         LED_128_Instance_addroundkey_out_36_,
         LED_128_Instance_addroundkey_out_37_,
         LED_128_Instance_addroundkey_out_38_,
         LED_128_Instance_addroundkey_out_48_,
         LED_128_Instance_addroundkey_out_49_,
         LED_128_Instance_addroundkey_out_50_,
         LED_128_Instance_addroundkey_out_51_,
         LED_128_Instance_addroundkey_out_52_,
         LED_128_Instance_addroundkey_out_53_,
         LED_128_Instance_addroundkey_out_54_, LED_128_Instance_n22,
         LED_128_Instance_MUX_current_roundkey_n10,
         LED_128_Instance_MUX_current_roundkey_n9,
         LED_128_Instance_MUX_current_roundkey_n8,
         LED_128_Instance_MUX_current_roundkey_n7,
         LED_128_Instance_MUX_addroundkey_out_n9,
         LED_128_Instance_MUX_addroundkey_out_n8,
         LED_128_Instance_MUX_addroundkey_out_n7,
         LED_128_Instance_SBox_Instance_0_n3,
         LED_128_Instance_SBox_Instance_0_n2,
         LED_128_Instance_SBox_Instance_0_n1,
         LED_128_Instance_SBox_Instance_0_L8,
         LED_128_Instance_SBox_Instance_0_L7,
         LED_128_Instance_SBox_Instance_0_T3,
         LED_128_Instance_SBox_Instance_0_T1,
         LED_128_Instance_SBox_Instance_0_Q7,
         LED_128_Instance_SBox_Instance_0_Q6,
         LED_128_Instance_SBox_Instance_0_L5,
         LED_128_Instance_SBox_Instance_0_T2,
         LED_128_Instance_SBox_Instance_0_L4,
         LED_128_Instance_SBox_Instance_0_Q3,
         LED_128_Instance_SBox_Instance_0_L3,
         LED_128_Instance_SBox_Instance_0_Q2,
         LED_128_Instance_SBox_Instance_0_T0,
         LED_128_Instance_SBox_Instance_0_L2,
         LED_128_Instance_SBox_Instance_0_L1,
         LED_128_Instance_SBox_Instance_0_L0,
         LED_128_Instance_SBox_Instance_1_n3,
         LED_128_Instance_SBox_Instance_1_n2,
         LED_128_Instance_SBox_Instance_1_n1,
         LED_128_Instance_SBox_Instance_1_L8,
         LED_128_Instance_SBox_Instance_1_L7,
         LED_128_Instance_SBox_Instance_1_T3,
         LED_128_Instance_SBox_Instance_1_T1,
         LED_128_Instance_SBox_Instance_1_Q7,
         LED_128_Instance_SBox_Instance_1_Q6,
         LED_128_Instance_SBox_Instance_1_L5,
         LED_128_Instance_SBox_Instance_1_T2,
         LED_128_Instance_SBox_Instance_1_L4,
         LED_128_Instance_SBox_Instance_1_Q3,
         LED_128_Instance_SBox_Instance_1_L3,
         LED_128_Instance_SBox_Instance_1_Q2,
         LED_128_Instance_SBox_Instance_1_T0,
         LED_128_Instance_SBox_Instance_1_L2,
         LED_128_Instance_SBox_Instance_1_L1,
         LED_128_Instance_SBox_Instance_1_L0,
         LED_128_Instance_SBox_Instance_2_n3,
         LED_128_Instance_SBox_Instance_2_n2,
         LED_128_Instance_SBox_Instance_2_n1,
         LED_128_Instance_SBox_Instance_2_L8,
         LED_128_Instance_SBox_Instance_2_L7,
         LED_128_Instance_SBox_Instance_2_T3,
         LED_128_Instance_SBox_Instance_2_T1,
         LED_128_Instance_SBox_Instance_2_Q7,
         LED_128_Instance_SBox_Instance_2_Q6,
         LED_128_Instance_SBox_Instance_2_L5,
         LED_128_Instance_SBox_Instance_2_T2,
         LED_128_Instance_SBox_Instance_2_L4,
         LED_128_Instance_SBox_Instance_2_Q3,
         LED_128_Instance_SBox_Instance_2_L3,
         LED_128_Instance_SBox_Instance_2_Q2,
         LED_128_Instance_SBox_Instance_2_T0,
         LED_128_Instance_SBox_Instance_2_L2,
         LED_128_Instance_SBox_Instance_2_L1,
         LED_128_Instance_SBox_Instance_2_L0,
         LED_128_Instance_SBox_Instance_3_n3,
         LED_128_Instance_SBox_Instance_3_n2,
         LED_128_Instance_SBox_Instance_3_n1,
         LED_128_Instance_SBox_Instance_3_L8,
         LED_128_Instance_SBox_Instance_3_L7,
         LED_128_Instance_SBox_Instance_3_T3,
         LED_128_Instance_SBox_Instance_3_T1,
         LED_128_Instance_SBox_Instance_3_Q7,
         LED_128_Instance_SBox_Instance_3_Q6,
         LED_128_Instance_SBox_Instance_3_L5,
         LED_128_Instance_SBox_Instance_3_T2,
         LED_128_Instance_SBox_Instance_3_L4,
         LED_128_Instance_SBox_Instance_3_Q3,
         LED_128_Instance_SBox_Instance_3_L3,
         LED_128_Instance_SBox_Instance_3_Q2,
         LED_128_Instance_SBox_Instance_3_T0,
         LED_128_Instance_SBox_Instance_3_L2,
         LED_128_Instance_SBox_Instance_3_L1,
         LED_128_Instance_SBox_Instance_3_L0,
         LED_128_Instance_SBox_Instance_4_n3,
         LED_128_Instance_SBox_Instance_4_n2,
         LED_128_Instance_SBox_Instance_4_n1,
         LED_128_Instance_SBox_Instance_4_L8,
         LED_128_Instance_SBox_Instance_4_L7,
         LED_128_Instance_SBox_Instance_4_T3,
         LED_128_Instance_SBox_Instance_4_T1,
         LED_128_Instance_SBox_Instance_4_Q7,
         LED_128_Instance_SBox_Instance_4_Q6,
         LED_128_Instance_SBox_Instance_4_L5,
         LED_128_Instance_SBox_Instance_4_T2,
         LED_128_Instance_SBox_Instance_4_L4,
         LED_128_Instance_SBox_Instance_4_Q3,
         LED_128_Instance_SBox_Instance_4_L3,
         LED_128_Instance_SBox_Instance_4_Q2,
         LED_128_Instance_SBox_Instance_4_T0,
         LED_128_Instance_SBox_Instance_4_L2,
         LED_128_Instance_SBox_Instance_4_L1,
         LED_128_Instance_SBox_Instance_4_L0,
         LED_128_Instance_SBox_Instance_5_n3,
         LED_128_Instance_SBox_Instance_5_n2,
         LED_128_Instance_SBox_Instance_5_n1,
         LED_128_Instance_SBox_Instance_5_L8,
         LED_128_Instance_SBox_Instance_5_L7,
         LED_128_Instance_SBox_Instance_5_T3,
         LED_128_Instance_SBox_Instance_5_T1,
         LED_128_Instance_SBox_Instance_5_Q7,
         LED_128_Instance_SBox_Instance_5_Q6,
         LED_128_Instance_SBox_Instance_5_L5,
         LED_128_Instance_SBox_Instance_5_T2,
         LED_128_Instance_SBox_Instance_5_L4,
         LED_128_Instance_SBox_Instance_5_Q3,
         LED_128_Instance_SBox_Instance_5_L3,
         LED_128_Instance_SBox_Instance_5_Q2,
         LED_128_Instance_SBox_Instance_5_T0,
         LED_128_Instance_SBox_Instance_5_L2,
         LED_128_Instance_SBox_Instance_5_L1,
         LED_128_Instance_SBox_Instance_5_L0,
         LED_128_Instance_SBox_Instance_6_n3,
         LED_128_Instance_SBox_Instance_6_n2,
         LED_128_Instance_SBox_Instance_6_n1,
         LED_128_Instance_SBox_Instance_6_L8,
         LED_128_Instance_SBox_Instance_6_L7,
         LED_128_Instance_SBox_Instance_6_T3,
         LED_128_Instance_SBox_Instance_6_T1,
         LED_128_Instance_SBox_Instance_6_Q7,
         LED_128_Instance_SBox_Instance_6_Q6,
         LED_128_Instance_SBox_Instance_6_L5,
         LED_128_Instance_SBox_Instance_6_T2,
         LED_128_Instance_SBox_Instance_6_L4,
         LED_128_Instance_SBox_Instance_6_Q3,
         LED_128_Instance_SBox_Instance_6_L3,
         LED_128_Instance_SBox_Instance_6_Q2,
         LED_128_Instance_SBox_Instance_6_T0,
         LED_128_Instance_SBox_Instance_6_L2,
         LED_128_Instance_SBox_Instance_6_L1,
         LED_128_Instance_SBox_Instance_6_L0,
         LED_128_Instance_SBox_Instance_7_n3,
         LED_128_Instance_SBox_Instance_7_n2,
         LED_128_Instance_SBox_Instance_7_n1,
         LED_128_Instance_SBox_Instance_7_L8,
         LED_128_Instance_SBox_Instance_7_L7,
         LED_128_Instance_SBox_Instance_7_T3,
         LED_128_Instance_SBox_Instance_7_T1,
         LED_128_Instance_SBox_Instance_7_Q7,
         LED_128_Instance_SBox_Instance_7_Q6,
         LED_128_Instance_SBox_Instance_7_L5,
         LED_128_Instance_SBox_Instance_7_T2,
         LED_128_Instance_SBox_Instance_7_L4,
         LED_128_Instance_SBox_Instance_7_Q3,
         LED_128_Instance_SBox_Instance_7_L3,
         LED_128_Instance_SBox_Instance_7_Q2,
         LED_128_Instance_SBox_Instance_7_T0,
         LED_128_Instance_SBox_Instance_7_L2,
         LED_128_Instance_SBox_Instance_7_L1,
         LED_128_Instance_SBox_Instance_7_L0,
         LED_128_Instance_SBox_Instance_8_n3,
         LED_128_Instance_SBox_Instance_8_n2,
         LED_128_Instance_SBox_Instance_8_n1,
         LED_128_Instance_SBox_Instance_8_L8,
         LED_128_Instance_SBox_Instance_8_L7,
         LED_128_Instance_SBox_Instance_8_T3,
         LED_128_Instance_SBox_Instance_8_T1,
         LED_128_Instance_SBox_Instance_8_Q7,
         LED_128_Instance_SBox_Instance_8_Q6,
         LED_128_Instance_SBox_Instance_8_L5,
         LED_128_Instance_SBox_Instance_8_T2,
         LED_128_Instance_SBox_Instance_8_L4,
         LED_128_Instance_SBox_Instance_8_Q3,
         LED_128_Instance_SBox_Instance_8_L3,
         LED_128_Instance_SBox_Instance_8_Q2,
         LED_128_Instance_SBox_Instance_8_T0,
         LED_128_Instance_SBox_Instance_8_L2,
         LED_128_Instance_SBox_Instance_8_L1,
         LED_128_Instance_SBox_Instance_8_L0,
         LED_128_Instance_SBox_Instance_9_n3,
         LED_128_Instance_SBox_Instance_9_n2,
         LED_128_Instance_SBox_Instance_9_n1,
         LED_128_Instance_SBox_Instance_9_L8,
         LED_128_Instance_SBox_Instance_9_L7,
         LED_128_Instance_SBox_Instance_9_T3,
         LED_128_Instance_SBox_Instance_9_T1,
         LED_128_Instance_SBox_Instance_9_Q7,
         LED_128_Instance_SBox_Instance_9_Q6,
         LED_128_Instance_SBox_Instance_9_L5,
         LED_128_Instance_SBox_Instance_9_T2,
         LED_128_Instance_SBox_Instance_9_L4,
         LED_128_Instance_SBox_Instance_9_Q3,
         LED_128_Instance_SBox_Instance_9_L3,
         LED_128_Instance_SBox_Instance_9_Q2,
         LED_128_Instance_SBox_Instance_9_T0,
         LED_128_Instance_SBox_Instance_9_L2,
         LED_128_Instance_SBox_Instance_9_L1,
         LED_128_Instance_SBox_Instance_9_L0,
         LED_128_Instance_SBox_Instance_10_n3,
         LED_128_Instance_SBox_Instance_10_n2,
         LED_128_Instance_SBox_Instance_10_n1,
         LED_128_Instance_SBox_Instance_10_L8,
         LED_128_Instance_SBox_Instance_10_L7,
         LED_128_Instance_SBox_Instance_10_T3,
         LED_128_Instance_SBox_Instance_10_T1,
         LED_128_Instance_SBox_Instance_10_Q7,
         LED_128_Instance_SBox_Instance_10_Q6,
         LED_128_Instance_SBox_Instance_10_L5,
         LED_128_Instance_SBox_Instance_10_T2,
         LED_128_Instance_SBox_Instance_10_L4,
         LED_128_Instance_SBox_Instance_10_Q3,
         LED_128_Instance_SBox_Instance_10_L3,
         LED_128_Instance_SBox_Instance_10_Q2,
         LED_128_Instance_SBox_Instance_10_T0,
         LED_128_Instance_SBox_Instance_10_L2,
         LED_128_Instance_SBox_Instance_10_L1,
         LED_128_Instance_SBox_Instance_10_L0,
         LED_128_Instance_SBox_Instance_11_n3,
         LED_128_Instance_SBox_Instance_11_n2,
         LED_128_Instance_SBox_Instance_11_n1,
         LED_128_Instance_SBox_Instance_11_L8,
         LED_128_Instance_SBox_Instance_11_L7,
         LED_128_Instance_SBox_Instance_11_T3,
         LED_128_Instance_SBox_Instance_11_T1,
         LED_128_Instance_SBox_Instance_11_Q7,
         LED_128_Instance_SBox_Instance_11_Q6,
         LED_128_Instance_SBox_Instance_11_L5,
         LED_128_Instance_SBox_Instance_11_T2,
         LED_128_Instance_SBox_Instance_11_L4,
         LED_128_Instance_SBox_Instance_11_Q3,
         LED_128_Instance_SBox_Instance_11_L3,
         LED_128_Instance_SBox_Instance_11_Q2,
         LED_128_Instance_SBox_Instance_11_T0,
         LED_128_Instance_SBox_Instance_11_L2,
         LED_128_Instance_SBox_Instance_11_L1,
         LED_128_Instance_SBox_Instance_11_L0,
         LED_128_Instance_SBox_Instance_12_n3,
         LED_128_Instance_SBox_Instance_12_n2,
         LED_128_Instance_SBox_Instance_12_n1,
         LED_128_Instance_SBox_Instance_12_L8,
         LED_128_Instance_SBox_Instance_12_L7,
         LED_128_Instance_SBox_Instance_12_T3,
         LED_128_Instance_SBox_Instance_12_T1,
         LED_128_Instance_SBox_Instance_12_Q7,
         LED_128_Instance_SBox_Instance_12_Q6,
         LED_128_Instance_SBox_Instance_12_L5,
         LED_128_Instance_SBox_Instance_12_T2,
         LED_128_Instance_SBox_Instance_12_L4,
         LED_128_Instance_SBox_Instance_12_Q3,
         LED_128_Instance_SBox_Instance_12_L3,
         LED_128_Instance_SBox_Instance_12_Q2,
         LED_128_Instance_SBox_Instance_12_T0,
         LED_128_Instance_SBox_Instance_12_L2,
         LED_128_Instance_SBox_Instance_12_L1,
         LED_128_Instance_SBox_Instance_12_L0,
         LED_128_Instance_SBox_Instance_13_n3,
         LED_128_Instance_SBox_Instance_13_n2,
         LED_128_Instance_SBox_Instance_13_n1,
         LED_128_Instance_SBox_Instance_13_L8,
         LED_128_Instance_SBox_Instance_13_L7,
         LED_128_Instance_SBox_Instance_13_T3,
         LED_128_Instance_SBox_Instance_13_T1,
         LED_128_Instance_SBox_Instance_13_Q7,
         LED_128_Instance_SBox_Instance_13_Q6,
         LED_128_Instance_SBox_Instance_13_L5,
         LED_128_Instance_SBox_Instance_13_T2,
         LED_128_Instance_SBox_Instance_13_L4,
         LED_128_Instance_SBox_Instance_13_Q3,
         LED_128_Instance_SBox_Instance_13_L3,
         LED_128_Instance_SBox_Instance_13_Q2,
         LED_128_Instance_SBox_Instance_13_T0,
         LED_128_Instance_SBox_Instance_13_L2,
         LED_128_Instance_SBox_Instance_13_L1,
         LED_128_Instance_SBox_Instance_13_L0,
         LED_128_Instance_SBox_Instance_14_n3,
         LED_128_Instance_SBox_Instance_14_n2,
         LED_128_Instance_SBox_Instance_14_n1,
         LED_128_Instance_SBox_Instance_14_L8,
         LED_128_Instance_SBox_Instance_14_L7,
         LED_128_Instance_SBox_Instance_14_T3,
         LED_128_Instance_SBox_Instance_14_T1,
         LED_128_Instance_SBox_Instance_14_Q7,
         LED_128_Instance_SBox_Instance_14_Q6,
         LED_128_Instance_SBox_Instance_14_L5,
         LED_128_Instance_SBox_Instance_14_T2,
         LED_128_Instance_SBox_Instance_14_L4,
         LED_128_Instance_SBox_Instance_14_Q3,
         LED_128_Instance_SBox_Instance_14_L3,
         LED_128_Instance_SBox_Instance_14_Q2,
         LED_128_Instance_SBox_Instance_14_T0,
         LED_128_Instance_SBox_Instance_14_L2,
         LED_128_Instance_SBox_Instance_14_L1,
         LED_128_Instance_SBox_Instance_14_L0,
         LED_128_Instance_SBox_Instance_15_n3,
         LED_128_Instance_SBox_Instance_15_n2,
         LED_128_Instance_SBox_Instance_15_n1,
         LED_128_Instance_SBox_Instance_15_L8,
         LED_128_Instance_SBox_Instance_15_L7,
         LED_128_Instance_SBox_Instance_15_T3,
         LED_128_Instance_SBox_Instance_15_T1,
         LED_128_Instance_SBox_Instance_15_Q7,
         LED_128_Instance_SBox_Instance_15_Q6,
         LED_128_Instance_SBox_Instance_15_L5,
         LED_128_Instance_SBox_Instance_15_T2,
         LED_128_Instance_SBox_Instance_15_L4,
         LED_128_Instance_SBox_Instance_15_Q3,
         LED_128_Instance_SBox_Instance_15_L3,
         LED_128_Instance_SBox_Instance_15_Q2,
         LED_128_Instance_SBox_Instance_15_T0,
         LED_128_Instance_SBox_Instance_15_L2,
         LED_128_Instance_SBox_Instance_15_L1,
         LED_128_Instance_SBox_Instance_15_L0,
         LED_128_Instance_MCS_Instance_0_n38,
         LED_128_Instance_MCS_Instance_0_n37,
         LED_128_Instance_MCS_Instance_0_n36,
         LED_128_Instance_MCS_Instance_0_n35,
         LED_128_Instance_MCS_Instance_0_n34,
         LED_128_Instance_MCS_Instance_0_n33,
         LED_128_Instance_MCS_Instance_0_n32,
         LED_128_Instance_MCS_Instance_0_n31,
         LED_128_Instance_MCS_Instance_0_n30,
         LED_128_Instance_MCS_Instance_0_n29,
         LED_128_Instance_MCS_Instance_0_n28,
         LED_128_Instance_MCS_Instance_0_n27,
         LED_128_Instance_MCS_Instance_0_n26,
         LED_128_Instance_MCS_Instance_0_n25,
         LED_128_Instance_MCS_Instance_0_n24,
         LED_128_Instance_MCS_Instance_0_n23,
         LED_128_Instance_MCS_Instance_0_n22,
         LED_128_Instance_MCS_Instance_0_n21,
         LED_128_Instance_MCS_Instance_0_n20,
         LED_128_Instance_MCS_Instance_0_n19,
         LED_128_Instance_MCS_Instance_0_n18,
         LED_128_Instance_MCS_Instance_0_n17,
         LED_128_Instance_MCS_Instance_0_n16,
         LED_128_Instance_MCS_Instance_0_n15,
         LED_128_Instance_MCS_Instance_0_n14,
         LED_128_Instance_MCS_Instance_0_n13,
         LED_128_Instance_MCS_Instance_0_n12,
         LED_128_Instance_MCS_Instance_0_n11,
         LED_128_Instance_MCS_Instance_0_n10,
         LED_128_Instance_MCS_Instance_0_n9,
         LED_128_Instance_MCS_Instance_0_n8,
         LED_128_Instance_MCS_Instance_0_n7,
         LED_128_Instance_MCS_Instance_0_n6,
         LED_128_Instance_MCS_Instance_0_n5,
         LED_128_Instance_MCS_Instance_0_n4,
         LED_128_Instance_MCS_Instance_0_n3,
         LED_128_Instance_MCS_Instance_0_n2,
         LED_128_Instance_MCS_Instance_0_n1,
         LED_128_Instance_MCS_Instance_1_n38,
         LED_128_Instance_MCS_Instance_1_n37,
         LED_128_Instance_MCS_Instance_1_n36,
         LED_128_Instance_MCS_Instance_1_n35,
         LED_128_Instance_MCS_Instance_1_n34,
         LED_128_Instance_MCS_Instance_1_n33,
         LED_128_Instance_MCS_Instance_1_n32,
         LED_128_Instance_MCS_Instance_1_n31,
         LED_128_Instance_MCS_Instance_1_n30,
         LED_128_Instance_MCS_Instance_1_n29,
         LED_128_Instance_MCS_Instance_1_n28,
         LED_128_Instance_MCS_Instance_1_n27,
         LED_128_Instance_MCS_Instance_1_n26,
         LED_128_Instance_MCS_Instance_1_n25,
         LED_128_Instance_MCS_Instance_1_n24,
         LED_128_Instance_MCS_Instance_1_n23,
         LED_128_Instance_MCS_Instance_1_n22,
         LED_128_Instance_MCS_Instance_1_n21,
         LED_128_Instance_MCS_Instance_1_n20,
         LED_128_Instance_MCS_Instance_1_n19,
         LED_128_Instance_MCS_Instance_1_n18,
         LED_128_Instance_MCS_Instance_1_n17,
         LED_128_Instance_MCS_Instance_1_n16,
         LED_128_Instance_MCS_Instance_1_n15,
         LED_128_Instance_MCS_Instance_1_n14,
         LED_128_Instance_MCS_Instance_1_n13,
         LED_128_Instance_MCS_Instance_1_n12,
         LED_128_Instance_MCS_Instance_1_n11,
         LED_128_Instance_MCS_Instance_1_n10,
         LED_128_Instance_MCS_Instance_1_n9,
         LED_128_Instance_MCS_Instance_1_n8,
         LED_128_Instance_MCS_Instance_1_n7,
         LED_128_Instance_MCS_Instance_1_n6,
         LED_128_Instance_MCS_Instance_1_n5,
         LED_128_Instance_MCS_Instance_1_n4,
         LED_128_Instance_MCS_Instance_1_n3,
         LED_128_Instance_MCS_Instance_1_n2,
         LED_128_Instance_MCS_Instance_1_n1,
         LED_128_Instance_MCS_Instance_2_n38,
         LED_128_Instance_MCS_Instance_2_n37,
         LED_128_Instance_MCS_Instance_2_n36,
         LED_128_Instance_MCS_Instance_2_n35,
         LED_128_Instance_MCS_Instance_2_n34,
         LED_128_Instance_MCS_Instance_2_n33,
         LED_128_Instance_MCS_Instance_2_n32,
         LED_128_Instance_MCS_Instance_2_n31,
         LED_128_Instance_MCS_Instance_2_n30,
         LED_128_Instance_MCS_Instance_2_n29,
         LED_128_Instance_MCS_Instance_2_n28,
         LED_128_Instance_MCS_Instance_2_n27,
         LED_128_Instance_MCS_Instance_2_n26,
         LED_128_Instance_MCS_Instance_2_n25,
         LED_128_Instance_MCS_Instance_2_n24,
         LED_128_Instance_MCS_Instance_2_n23,
         LED_128_Instance_MCS_Instance_2_n22,
         LED_128_Instance_MCS_Instance_2_n21,
         LED_128_Instance_MCS_Instance_2_n20,
         LED_128_Instance_MCS_Instance_2_n19,
         LED_128_Instance_MCS_Instance_2_n18,
         LED_128_Instance_MCS_Instance_2_n17,
         LED_128_Instance_MCS_Instance_2_n16,
         LED_128_Instance_MCS_Instance_2_n15,
         LED_128_Instance_MCS_Instance_2_n14,
         LED_128_Instance_MCS_Instance_2_n13,
         LED_128_Instance_MCS_Instance_2_n12,
         LED_128_Instance_MCS_Instance_2_n11,
         LED_128_Instance_MCS_Instance_2_n10,
         LED_128_Instance_MCS_Instance_2_n9,
         LED_128_Instance_MCS_Instance_2_n8,
         LED_128_Instance_MCS_Instance_2_n7,
         LED_128_Instance_MCS_Instance_2_n6,
         LED_128_Instance_MCS_Instance_2_n5,
         LED_128_Instance_MCS_Instance_2_n4,
         LED_128_Instance_MCS_Instance_2_n3,
         LED_128_Instance_MCS_Instance_2_n2,
         LED_128_Instance_MCS_Instance_2_n1,
         LED_128_Instance_MCS_Instance_3_n38,
         LED_128_Instance_MCS_Instance_3_n37,
         LED_128_Instance_MCS_Instance_3_n36,
         LED_128_Instance_MCS_Instance_3_n35,
         LED_128_Instance_MCS_Instance_3_n34,
         LED_128_Instance_MCS_Instance_3_n33,
         LED_128_Instance_MCS_Instance_3_n32,
         LED_128_Instance_MCS_Instance_3_n31,
         LED_128_Instance_MCS_Instance_3_n30,
         LED_128_Instance_MCS_Instance_3_n29,
         LED_128_Instance_MCS_Instance_3_n28,
         LED_128_Instance_MCS_Instance_3_n27,
         LED_128_Instance_MCS_Instance_3_n26,
         LED_128_Instance_MCS_Instance_3_n25,
         LED_128_Instance_MCS_Instance_3_n24,
         LED_128_Instance_MCS_Instance_3_n23,
         LED_128_Instance_MCS_Instance_3_n22,
         LED_128_Instance_MCS_Instance_3_n21,
         LED_128_Instance_MCS_Instance_3_n20,
         LED_128_Instance_MCS_Instance_3_n19,
         LED_128_Instance_MCS_Instance_3_n18,
         LED_128_Instance_MCS_Instance_3_n17,
         LED_128_Instance_MCS_Instance_3_n16,
         LED_128_Instance_MCS_Instance_3_n15,
         LED_128_Instance_MCS_Instance_3_n14,
         LED_128_Instance_MCS_Instance_3_n13,
         LED_128_Instance_MCS_Instance_3_n12,
         LED_128_Instance_MCS_Instance_3_n11,
         LED_128_Instance_MCS_Instance_3_n10,
         LED_128_Instance_MCS_Instance_3_n9,
         LED_128_Instance_MCS_Instance_3_n8,
         LED_128_Instance_MCS_Instance_3_n7,
         LED_128_Instance_MCS_Instance_3_n6,
         LED_128_Instance_MCS_Instance_3_n5,
         LED_128_Instance_MCS_Instance_3_n4,
         LED_128_Instance_MCS_Instance_3_n3,
         LED_128_Instance_MCS_Instance_3_n2,
         LED_128_Instance_MCS_Instance_3_n1, LED_128_Instance_ks_reg_0__Q,
         LED_128_Instance_cipherstate_reg_0__QN,
         LED_128_Instance_cipherstate_reg_1__QN,
         LED_128_Instance_cipherstate_reg_2__QN,
         LED_128_Instance_cipherstate_reg_3__QN,
         LED_128_Instance_cipherstate_reg_4__QN,
         LED_128_Instance_cipherstate_reg_5__QN,
         LED_128_Instance_cipherstate_reg_6__QN,
         LED_128_Instance_cipherstate_reg_7__QN,
         LED_128_Instance_cipherstate_reg_8__QN,
         LED_128_Instance_cipherstate_reg_9__QN,
         LED_128_Instance_cipherstate_reg_10__QN,
         LED_128_Instance_cipherstate_reg_11__QN,
         LED_128_Instance_cipherstate_reg_12__QN,
         LED_128_Instance_cipherstate_reg_13__QN,
         LED_128_Instance_cipherstate_reg_14__QN,
         LED_128_Instance_cipherstate_reg_15__QN,
         LED_128_Instance_cipherstate_reg_16__QN,
         LED_128_Instance_cipherstate_reg_17__QN,
         LED_128_Instance_cipherstate_reg_18__QN,
         LED_128_Instance_cipherstate_reg_19__QN,
         LED_128_Instance_cipherstate_reg_20__QN,
         LED_128_Instance_cipherstate_reg_21__QN,
         LED_128_Instance_cipherstate_reg_22__QN,
         LED_128_Instance_cipherstate_reg_23__QN,
         LED_128_Instance_cipherstate_reg_24__QN,
         LED_128_Instance_cipherstate_reg_25__QN,
         LED_128_Instance_cipherstate_reg_26__QN,
         LED_128_Instance_cipherstate_reg_27__QN,
         LED_128_Instance_cipherstate_reg_28__QN,
         LED_128_Instance_cipherstate_reg_29__QN,
         LED_128_Instance_cipherstate_reg_30__QN,
         LED_128_Instance_cipherstate_reg_31__QN,
         LED_128_Instance_cipherstate_reg_32__QN,
         LED_128_Instance_cipherstate_reg_33__QN,
         LED_128_Instance_cipherstate_reg_34__QN,
         LED_128_Instance_cipherstate_reg_35__QN,
         LED_128_Instance_cipherstate_reg_36__QN,
         LED_128_Instance_cipherstate_reg_37__QN,
         LED_128_Instance_cipherstate_reg_38__QN,
         LED_128_Instance_cipherstate_reg_39__QN,
         LED_128_Instance_cipherstate_reg_40__QN,
         LED_128_Instance_cipherstate_reg_41__QN,
         LED_128_Instance_cipherstate_reg_42__QN,
         LED_128_Instance_cipherstate_reg_43__QN,
         LED_128_Instance_cipherstate_reg_44__QN,
         LED_128_Instance_cipherstate_reg_45__QN,
         LED_128_Instance_cipherstate_reg_46__QN,
         LED_128_Instance_cipherstate_reg_47__QN,
         LED_128_Instance_cipherstate_reg_48__QN,
         LED_128_Instance_cipherstate_reg_49__QN,
         LED_128_Instance_cipherstate_reg_50__QN,
         LED_128_Instance_cipherstate_reg_51__QN,
         LED_128_Instance_cipherstate_reg_52__QN,
         LED_128_Instance_cipherstate_reg_53__QN,
         LED_128_Instance_cipherstate_reg_54__QN,
         LED_128_Instance_cipherstate_reg_55__QN,
         LED_128_Instance_cipherstate_reg_56__QN,
         LED_128_Instance_cipherstate_reg_57__QN,
         LED_128_Instance_cipherstate_reg_58__QN,
         LED_128_Instance_cipherstate_reg_59__QN,
         LED_128_Instance_cipherstate_reg_60__QN,
         LED_128_Instance_cipherstate_reg_61__QN,
         LED_128_Instance_cipherstate_reg_62__QN,
         LED_128_Instance_cipherstate_reg_63__QN, internal_done_reg_QN;
  wire   [5:0] roundconstant;
  (* AGEMA = "layer" *) wire LED_128_Instance_MUX_state0_n11;
  (* AGEMA = "layer" *) wire LED_128_Instance_MUX_state0_n10;
  (* AGEMA = "layer" *) wire LED_128_Instance_MUX_state0_n9;
  (* AGEMA = "layer" *) wire LED_128_Instance_MUX_state0_n8;
  (* AGEMA = "layer" *) wire   [63:0] LED_128_Instance_subcells_out;
  (* AGEMA = "layer" *) wire   [63:0] LED_128_Instance_addconst_out;
  (* AGEMA = "layer" *) wire   [63:0] LED_128_Instance_addroundkey_tmp;
  wire   [63:0] LED_128_Instance_current_roundkey;
  wire   [63:0] LED_128_Instance_state1;
  wire   [63:0] LED_128_Instance_state0;
  wire   [63:0] LED_128_Instance_mixcolumns_out;

  NOR2_X1 U16 ( .A1(roundconstant[4]), .A2(roundconstant[1]), .ZN(n14) );
  NAND2_X1 U17 ( .A1(roundconstant[0]), .A2(n14), .ZN(n16) );
  NOR2_X1 U18 ( .A1(roundconstant[5]), .A2(n16), .ZN(n17) );
  NAND2_X1 U19 ( .A1(roundconstant[3]), .A2(n17), .ZN(n18) );
  NOR2_X1 U20 ( .A1(roundconstant[2]), .A2(n18), .ZN(n19) );
  NOR2_X1 U21 ( .A1(OUT_done), .A2(n19), .ZN(n20) );
  NOR2_X1 U22 ( .A1(IN_reset), .A2(n20), .ZN(n15) );
  NAND2_X1 LED_128_Instance_U30 ( .A1(LED_128_Instance_n33), .A2(
        LED_128_Instance_n32), .ZN(LED_128_Instance_n34) );
  XNOR2_X1 LED_128_Instance_U29 ( .A(LED_128_Instance_n25), .B(
        LED_128_Instance_n23), .ZN(LED_128_Instance_n32) );
  XOR2_X1 LED_128_Instance_U28 ( .A(LED_128_Instance_n4), .B(
        LED_128_Instance_n26), .Z(LED_128_Instance_n23) );
  NAND2_X1 LED_128_Instance_U27 ( .A1(LED_128_Instance_n21), .A2(
        LED_128_Instance_n20), .ZN(LED_128_Instance_n33) );
  NAND2_X1 LED_128_Instance_U26 ( .A1(LED_128_Instance_n19), .A2(
        LED_128_Instance_n18), .ZN(LED_128_Instance_n20) );
  NOR2_X1 LED_128_Instance_U25 ( .A1(LED_128_Instance_n24), .A2(
        LED_128_Instance_n1), .ZN(LED_128_Instance_n18) );
  NOR2_X1 LED_128_Instance_U24 ( .A1(LED_128_Instance_n8), .A2(
        LED_128_Instance_n4), .ZN(LED_128_Instance_n19) );
  NAND2_X1 LED_128_Instance_U23 ( .A1(LED_128_Instance_n1), .A2(
        LED_128_Instance_n17), .ZN(LED_128_Instance_n21) );
  AND2_X1 LED_128_Instance_U22 ( .A1(LED_128_Instance_n8), .A2(
        LED_128_Instance_n4), .ZN(LED_128_Instance_n17) );
  NAND2_X1 LED_128_Instance_U21 ( .A1(LED_128_Instance_n29), .A2(
        LED_128_Instance_n14), .ZN(LED_128_Instance_n15) );
  NOR2_X1 LED_128_Instance_U20 ( .A1(LED_128_Instance_n6), .A2(
        LED_128_Instance_n13), .ZN(LED_128_Instance_n14) );
  NAND2_X1 LED_128_Instance_U19 ( .A1(LED_128_Instance_n5), .A2(
        roundconstant[3]), .ZN(LED_128_Instance_n13) );
  NAND2_X1 LED_128_Instance_U18 ( .A1(LED_128_Instance_n28), .A2(
        LED_128_Instance_n27), .ZN(LED_128_Instance_n16) );
  NOR2_X1 LED_128_Instance_U17 ( .A1(LED_128_Instance_n28), .A2(IN_reset), 
        .ZN(LED_128_Instance_N9) );
  NOR2_X1 LED_128_Instance_U16 ( .A1(IN_reset), .A2(LED_128_Instance_n30), 
        .ZN(LED_128_Instance_N8) );
  NOR2_X1 LED_128_Instance_U15 ( .A1(IN_reset), .A2(LED_128_Instance_n5), .ZN(
        LED_128_Instance_N7) );
  NOR2_X1 LED_128_Instance_U14 ( .A1(IN_reset), .A2(LED_128_Instance_n29), 
        .ZN(LED_128_Instance_N6) );
  NOR2_X1 LED_128_Instance_U13 ( .A1(IN_reset), .A2(LED_128_Instance_n6), .ZN(
        LED_128_Instance_N5) );
  NOR2_X1 LED_128_Instance_U12 ( .A1(LED_128_Instance_n1), .A2(IN_reset), .ZN(
        LED_128_Instance_N13) );
  NOR2_X1 LED_128_Instance_U11 ( .A1(LED_128_Instance_n8), .A2(IN_reset), .ZN(
        LED_128_Instance_N12) );
  NOR2_X1 LED_128_Instance_U10 ( .A1(LED_128_Instance_n4), .A2(IN_reset), .ZN(
        LED_128_Instance_N11) );
  NOR2_X1 LED_128_Instance_U9 ( .A1(LED_128_Instance_n2), .A2(IN_reset), .ZN(
        LED_128_Instance_N10) );
  OR2_X1 LED_128_Instance_U8 ( .A1(LED_128_Instance_n2), .A2(
        LED_128_Instance_n21), .ZN(LED_128_Instance_n11) );
  NAND2_X1 LED_128_Instance_U7 ( .A1(LED_128_Instance_n34), .A2(
        LED_128_Instance_n11), .ZN(LED_128_Instance_n31) );
  NOR2_X1 LED_128_Instance_U6 ( .A1(LED_128_Instance_n16), .A2(
        LED_128_Instance_n15), .ZN(LED_128_Instance_n22) );
  INV_X1 LED_128_Instance_U5 ( .A(LED_128_Instance_n11), .ZN(
        LED_128_Instance_n12) );
  OR2_X1 LED_128_Instance_U4 ( .A1(IN_reset), .A2(LED_128_Instance_n10), .ZN(
        LED_128_Instance_N4) );
  XNOR2_X1 LED_128_Instance_U3 ( .A(LED_128_Instance_n28), .B(
        LED_128_Instance_n27), .ZN(LED_128_Instance_n10) );
  INV_X1 LED_128_Instance_MUX_state0_U4 ( .A(LED_128_Instance_n22), .ZN(
        LED_128_Instance_MUX_state0_n11) );
  INV_X1 LED_128_Instance_MUX_state0_U3 ( .A(LED_128_Instance_MUX_state0_n11), 
        .ZN(LED_128_Instance_MUX_state0_n8) );
  INV_X1 LED_128_Instance_MUX_state0_U2 ( .A(LED_128_Instance_MUX_state0_n11), 
        .ZN(LED_128_Instance_MUX_state0_n10) );
  INV_X1 LED_128_Instance_MUX_state0_U1 ( .A(LED_128_Instance_MUX_state0_n11), 
        .ZN(LED_128_Instance_MUX_state0_n9) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_0_U1 ( .A(
        LED_128_Instance_mixcolumns_out[0]), .B(
        LED_128_Instance_addroundkey_out_0_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[0]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_1_U1 ( .A(
        LED_128_Instance_mixcolumns_out[1]), .B(
        LED_128_Instance_addroundkey_out_1_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[1]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_2_U1 ( .A(
        LED_128_Instance_mixcolumns_out[2]), .B(
        LED_128_Instance_addroundkey_out_2_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[2]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_3_U1 ( .A(
        LED_128_Instance_mixcolumns_out[3]), .B(
        LED_128_Instance_addroundkey_out_3_), .S(
        LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[3]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_4_U1 ( .A(
        LED_128_Instance_mixcolumns_out[4]), .B(
        LED_128_Instance_addroundkey_out_4_), .S(
        LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[4]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_5_U1 ( .A(
        LED_128_Instance_mixcolumns_out[5]), .B(
        LED_128_Instance_addroundkey_out_5_), .S(
        LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[5]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_6_U1 ( .A(
        LED_128_Instance_mixcolumns_out[6]), .B(
        LED_128_Instance_addroundkey_out_6_), .S(
        LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[6]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_7_U1 ( .A(
        LED_128_Instance_mixcolumns_out[7]), .B(
        LED_128_Instance_addconst_out[7]), .S(LED_128_Instance_MUX_state0_n10), 
        .Z(LED_128_Instance_state0[7]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_8_U1 ( .A(
        LED_128_Instance_mixcolumns_out[8]), .B(
        LED_128_Instance_addconst_out[8]), .S(LED_128_Instance_MUX_state0_n10), 
        .Z(LED_128_Instance_state0[8]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_9_U1 ( .A(
        LED_128_Instance_mixcolumns_out[9]), .B(
        LED_128_Instance_addconst_out[9]), .S(LED_128_Instance_MUX_state0_n10), 
        .Z(LED_128_Instance_state0[9]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_10_U1 ( .A(
        LED_128_Instance_mixcolumns_out[10]), .B(
        LED_128_Instance_addconst_out[10]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[10]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_11_U1 ( .A(
        LED_128_Instance_mixcolumns_out[11]), .B(
        LED_128_Instance_addconst_out[11]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[11]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_12_U1 ( .A(
        LED_128_Instance_mixcolumns_out[12]), .B(
        LED_128_Instance_addconst_out[12]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[12]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_13_U1 ( .A(
        LED_128_Instance_mixcolumns_out[13]), .B(
        LED_128_Instance_addconst_out[13]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[13]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_14_U1 ( .A(
        LED_128_Instance_mixcolumns_out[14]), .B(
        LED_128_Instance_addconst_out[14]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[14]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_15_U1 ( .A(
        LED_128_Instance_mixcolumns_out[15]), .B(
        LED_128_Instance_addconst_out[15]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[15]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_16_U1 ( .A(
        LED_128_Instance_mixcolumns_out[16]), .B(
        LED_128_Instance_addroundkey_out_16_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[16]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_17_U1 ( .A(
        LED_128_Instance_mixcolumns_out[17]), .B(
        LED_128_Instance_addroundkey_out_17_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[17]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_18_U1 ( .A(
        LED_128_Instance_mixcolumns_out[18]), .B(
        LED_128_Instance_addroundkey_out_18_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[18]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_19_U1 ( .A(
        LED_128_Instance_mixcolumns_out[19]), .B(
        LED_128_Instance_addroundkey_out_19_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[19]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_20_U1 ( .A(
        LED_128_Instance_mixcolumns_out[20]), .B(
        LED_128_Instance_addroundkey_out_20_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[20]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_21_U1 ( .A(
        LED_128_Instance_mixcolumns_out[21]), .B(
        LED_128_Instance_addroundkey_out_21_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[21]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_22_U1 ( .A(
        LED_128_Instance_mixcolumns_out[22]), .B(
        LED_128_Instance_addroundkey_out_22_), .S(
        LED_128_Instance_MUX_state0_n9), .Z(LED_128_Instance_state0[22]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_23_U1 ( .A(
        LED_128_Instance_mixcolumns_out[23]), .B(
        LED_128_Instance_addconst_out[23]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[23]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_24_U1 ( .A(
        LED_128_Instance_mixcolumns_out[24]), .B(
        LED_128_Instance_addconst_out[24]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[24]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_25_U1 ( .A(
        LED_128_Instance_mixcolumns_out[25]), .B(
        LED_128_Instance_addconst_out[25]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[25]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_26_U1 ( .A(
        LED_128_Instance_mixcolumns_out[26]), .B(
        LED_128_Instance_addconst_out[26]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[26]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_27_U1 ( .A(
        LED_128_Instance_mixcolumns_out[27]), .B(
        LED_128_Instance_addconst_out[27]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[27]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_28_U1 ( .A(
        LED_128_Instance_mixcolumns_out[28]), .B(
        LED_128_Instance_addconst_out[28]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[28]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_29_U1 ( .A(
        LED_128_Instance_mixcolumns_out[29]), .B(
        LED_128_Instance_addconst_out[29]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[29]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_30_U1 ( .A(
        LED_128_Instance_mixcolumns_out[30]), .B(
        LED_128_Instance_addconst_out[30]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[30]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_31_U1 ( .A(
        LED_128_Instance_mixcolumns_out[31]), .B(
        LED_128_Instance_addconst_out[31]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[31]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_32_U1 ( .A(
        LED_128_Instance_mixcolumns_out[32]), .B(
        LED_128_Instance_addroundkey_out_32_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[32]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_33_U1 ( .A(
        LED_128_Instance_mixcolumns_out[33]), .B(
        LED_128_Instance_addroundkey_out_33_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[33]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_34_U1 ( .A(
        LED_128_Instance_mixcolumns_out[34]), .B(
        LED_128_Instance_addroundkey_out_34_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[34]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_35_U1 ( .A(
        LED_128_Instance_mixcolumns_out[35]), .B(
        LED_128_Instance_addroundkey_out_35_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[35]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_36_U1 ( .A(
        LED_128_Instance_mixcolumns_out[36]), .B(
        LED_128_Instance_addroundkey_out_36_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[36]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_37_U1 ( .A(
        LED_128_Instance_mixcolumns_out[37]), .B(
        LED_128_Instance_addroundkey_out_37_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[37]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_38_U1 ( .A(
        LED_128_Instance_mixcolumns_out[38]), .B(
        LED_128_Instance_addroundkey_out_38_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[38]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_39_U1 ( .A(
        LED_128_Instance_mixcolumns_out[39]), .B(
        LED_128_Instance_addconst_out[39]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[39]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_40_U1 ( .A(
        LED_128_Instance_mixcolumns_out[40]), .B(
        LED_128_Instance_addconst_out[40]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[40]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_41_U1 ( .A(
        LED_128_Instance_mixcolumns_out[41]), .B(
        LED_128_Instance_addconst_out[41]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[41]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_42_U1 ( .A(
        LED_128_Instance_mixcolumns_out[42]), .B(
        LED_128_Instance_addconst_out[42]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[42]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_43_U1 ( .A(
        LED_128_Instance_mixcolumns_out[43]), .B(
        LED_128_Instance_addconst_out[43]), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[43]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_44_U1 ( .A(
        LED_128_Instance_mixcolumns_out[44]), .B(
        LED_128_Instance_addconst_out[44]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[44]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_45_U1 ( .A(
        LED_128_Instance_mixcolumns_out[45]), .B(
        LED_128_Instance_addconst_out[45]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[45]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_46_U1 ( .A(
        LED_128_Instance_mixcolumns_out[46]), .B(
        LED_128_Instance_addconst_out[46]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[46]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_47_U1 ( .A(
        LED_128_Instance_mixcolumns_out[47]), .B(
        LED_128_Instance_addconst_out[47]), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[47]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_48_U1 ( .A(
        LED_128_Instance_mixcolumns_out[48]), .B(
        LED_128_Instance_addroundkey_out_48_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[48]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_49_U1 ( .A(
        LED_128_Instance_mixcolumns_out[49]), .B(
        LED_128_Instance_addroundkey_out_49_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[49]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_50_U1 ( .A(
        LED_128_Instance_mixcolumns_out[50]), .B(
        LED_128_Instance_addroundkey_out_50_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[50]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_51_U1 ( .A(
        LED_128_Instance_mixcolumns_out[51]), .B(
        LED_128_Instance_addroundkey_out_51_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[51]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_52_U1 ( .A(
        LED_128_Instance_mixcolumns_out[52]), .B(
        LED_128_Instance_addroundkey_out_52_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[52]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_53_U1 ( .A(
        LED_128_Instance_mixcolumns_out[53]), .B(
        LED_128_Instance_addroundkey_out_53_), .S(LED_128_Instance_n22), .Z(
        LED_128_Instance_state0[53]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_54_U1 ( .A(
        LED_128_Instance_mixcolumns_out[54]), .B(
        LED_128_Instance_addroundkey_out_54_), .S(
        LED_128_Instance_MUX_state0_n8), .Z(LED_128_Instance_state0[54]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_55_U1 ( .A(
        LED_128_Instance_mixcolumns_out[55]), .B(
        LED_128_Instance_addconst_out[55]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[55]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_56_U1 ( .A(
        LED_128_Instance_mixcolumns_out[56]), .B(
        LED_128_Instance_addconst_out[56]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[56]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_57_U1 ( .A(
        LED_128_Instance_mixcolumns_out[57]), .B(
        LED_128_Instance_addconst_out[57]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[57]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_58_U1 ( .A(
        LED_128_Instance_mixcolumns_out[58]), .B(
        LED_128_Instance_addconst_out[58]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[58]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_59_U1 ( .A(
        LED_128_Instance_mixcolumns_out[59]), .B(
        LED_128_Instance_addconst_out[59]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[59]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_60_U1 ( .A(
        LED_128_Instance_mixcolumns_out[60]), .B(
        LED_128_Instance_addconst_out[60]), .S(LED_128_Instance_MUX_state0_n9), 
        .Z(LED_128_Instance_state0[60]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_61_U1 ( .A(
        LED_128_Instance_mixcolumns_out[61]), .B(
        LED_128_Instance_addconst_out[61]), .S(LED_128_Instance_MUX_state0_n10), .Z(LED_128_Instance_state0[61]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_62_U1 ( .A(
        LED_128_Instance_mixcolumns_out[62]), .B(
        LED_128_Instance_addconst_out[62]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[62]) );
  MUX2_X1 LED_128_Instance_MUX_state0_mux_inst_63_U1 ( .A(
        LED_128_Instance_mixcolumns_out[63]), .B(
        LED_128_Instance_addconst_out[63]), .S(LED_128_Instance_MUX_state0_n8), 
        .Z(LED_128_Instance_state0[63]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_0_U1 ( .A(
        LED_128_Instance_state0[0]), .B(IN_plaintext[0]), .S(IN_reset), .Z(
        LED_128_Instance_state1[0]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_1_U1 ( .A(
        LED_128_Instance_state0[1]), .B(IN_plaintext[1]), .S(IN_reset), .Z(
        LED_128_Instance_state1[1]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_2_U1 ( .A(
        LED_128_Instance_state0[2]), .B(IN_plaintext[2]), .S(IN_reset), .Z(
        LED_128_Instance_state1[2]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_3_U1 ( .A(
        LED_128_Instance_state0[3]), .B(IN_plaintext[3]), .S(IN_reset), .Z(
        LED_128_Instance_state1[3]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_4_U1 ( .A(
        LED_128_Instance_state0[4]), .B(IN_plaintext[4]), .S(IN_reset), .Z(
        LED_128_Instance_state1[4]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_5_U1 ( .A(
        LED_128_Instance_state0[5]), .B(IN_plaintext[5]), .S(IN_reset), .Z(
        LED_128_Instance_state1[5]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_6_U1 ( .A(
        LED_128_Instance_state0[6]), .B(IN_plaintext[6]), .S(IN_reset), .Z(
        LED_128_Instance_state1[6]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_7_U1 ( .A(
        LED_128_Instance_state0[7]), .B(IN_plaintext[7]), .S(IN_reset), .Z(
        LED_128_Instance_state1[7]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_8_U1 ( .A(
        LED_128_Instance_state0[8]), .B(IN_plaintext[8]), .S(IN_reset), .Z(
        LED_128_Instance_state1[8]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_9_U1 ( .A(
        LED_128_Instance_state0[9]), .B(IN_plaintext[9]), .S(IN_reset), .Z(
        LED_128_Instance_state1[9]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_10_U1 ( .A(
        LED_128_Instance_state0[10]), .B(IN_plaintext[10]), .S(IN_reset), .Z(
        LED_128_Instance_state1[10]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_11_U1 ( .A(
        LED_128_Instance_state0[11]), .B(IN_plaintext[11]), .S(IN_reset), .Z(
        LED_128_Instance_state1[11]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_12_U1 ( .A(
        LED_128_Instance_state0[12]), .B(IN_plaintext[12]), .S(IN_reset), .Z(
        LED_128_Instance_state1[12]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_13_U1 ( .A(
        LED_128_Instance_state0[13]), .B(IN_plaintext[13]), .S(IN_reset), .Z(
        LED_128_Instance_state1[13]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_14_U1 ( .A(
        LED_128_Instance_state0[14]), .B(IN_plaintext[14]), .S(IN_reset), .Z(
        LED_128_Instance_state1[14]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_15_U1 ( .A(
        LED_128_Instance_state0[15]), .B(IN_plaintext[15]), .S(IN_reset), .Z(
        LED_128_Instance_state1[15]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_16_U1 ( .A(
        LED_128_Instance_state0[16]), .B(IN_plaintext[16]), .S(IN_reset), .Z(
        LED_128_Instance_state1[16]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_17_U1 ( .A(
        LED_128_Instance_state0[17]), .B(IN_plaintext[17]), .S(IN_reset), .Z(
        LED_128_Instance_state1[17]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_18_U1 ( .A(
        LED_128_Instance_state0[18]), .B(IN_plaintext[18]), .S(IN_reset), .Z(
        LED_128_Instance_state1[18]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_19_U1 ( .A(
        LED_128_Instance_state0[19]), .B(IN_plaintext[19]), .S(IN_reset), .Z(
        LED_128_Instance_state1[19]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_20_U1 ( .A(
        LED_128_Instance_state0[20]), .B(IN_plaintext[20]), .S(IN_reset), .Z(
        LED_128_Instance_state1[20]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_21_U1 ( .A(
        LED_128_Instance_state0[21]), .B(IN_plaintext[21]), .S(IN_reset), .Z(
        LED_128_Instance_state1[21]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_22_U1 ( .A(
        LED_128_Instance_state0[22]), .B(IN_plaintext[22]), .S(IN_reset), .Z(
        LED_128_Instance_state1[22]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_23_U1 ( .A(
        LED_128_Instance_state0[23]), .B(IN_plaintext[23]), .S(IN_reset), .Z(
        LED_128_Instance_state1[23]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_24_U1 ( .A(
        LED_128_Instance_state0[24]), .B(IN_plaintext[24]), .S(IN_reset), .Z(
        LED_128_Instance_state1[24]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_25_U1 ( .A(
        LED_128_Instance_state0[25]), .B(IN_plaintext[25]), .S(IN_reset), .Z(
        LED_128_Instance_state1[25]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_26_U1 ( .A(
        LED_128_Instance_state0[26]), .B(IN_plaintext[26]), .S(IN_reset), .Z(
        LED_128_Instance_state1[26]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_27_U1 ( .A(
        LED_128_Instance_state0[27]), .B(IN_plaintext[27]), .S(IN_reset), .Z(
        LED_128_Instance_state1[27]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_28_U1 ( .A(
        LED_128_Instance_state0[28]), .B(IN_plaintext[28]), .S(IN_reset), .Z(
        LED_128_Instance_state1[28]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_29_U1 ( .A(
        LED_128_Instance_state0[29]), .B(IN_plaintext[29]), .S(IN_reset), .Z(
        LED_128_Instance_state1[29]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_30_U1 ( .A(
        LED_128_Instance_state0[30]), .B(IN_plaintext[30]), .S(IN_reset), .Z(
        LED_128_Instance_state1[30]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_31_U1 ( .A(
        LED_128_Instance_state0[31]), .B(IN_plaintext[31]), .S(IN_reset), .Z(
        LED_128_Instance_state1[31]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_32_U1 ( .A(
        LED_128_Instance_state0[32]), .B(IN_plaintext[32]), .S(IN_reset), .Z(
        LED_128_Instance_state1[32]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_33_U1 ( .A(
        LED_128_Instance_state0[33]), .B(IN_plaintext[33]), .S(IN_reset), .Z(
        LED_128_Instance_state1[33]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_34_U1 ( .A(
        LED_128_Instance_state0[34]), .B(IN_plaintext[34]), .S(IN_reset), .Z(
        LED_128_Instance_state1[34]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_35_U1 ( .A(
        LED_128_Instance_state0[35]), .B(IN_plaintext[35]), .S(IN_reset), .Z(
        LED_128_Instance_state1[35]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_36_U1 ( .A(
        LED_128_Instance_state0[36]), .B(IN_plaintext[36]), .S(IN_reset), .Z(
        LED_128_Instance_state1[36]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_37_U1 ( .A(
        LED_128_Instance_state0[37]), .B(IN_plaintext[37]), .S(IN_reset), .Z(
        LED_128_Instance_state1[37]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_38_U1 ( .A(
        LED_128_Instance_state0[38]), .B(IN_plaintext[38]), .S(IN_reset), .Z(
        LED_128_Instance_state1[38]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_39_U1 ( .A(
        LED_128_Instance_state0[39]), .B(IN_plaintext[39]), .S(IN_reset), .Z(
        LED_128_Instance_state1[39]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_40_U1 ( .A(
        LED_128_Instance_state0[40]), .B(IN_plaintext[40]), .S(IN_reset), .Z(
        LED_128_Instance_state1[40]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_41_U1 ( .A(
        LED_128_Instance_state0[41]), .B(IN_plaintext[41]), .S(IN_reset), .Z(
        LED_128_Instance_state1[41]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_42_U1 ( .A(
        LED_128_Instance_state0[42]), .B(IN_plaintext[42]), .S(IN_reset), .Z(
        LED_128_Instance_state1[42]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_43_U1 ( .A(
        LED_128_Instance_state0[43]), .B(IN_plaintext[43]), .S(IN_reset), .Z(
        LED_128_Instance_state1[43]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_44_U1 ( .A(
        LED_128_Instance_state0[44]), .B(IN_plaintext[44]), .S(IN_reset), .Z(
        LED_128_Instance_state1[44]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_45_U1 ( .A(
        LED_128_Instance_state0[45]), .B(IN_plaintext[45]), .S(IN_reset), .Z(
        LED_128_Instance_state1[45]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_46_U1 ( .A(
        LED_128_Instance_state0[46]), .B(IN_plaintext[46]), .S(IN_reset), .Z(
        LED_128_Instance_state1[46]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_47_U1 ( .A(
        LED_128_Instance_state0[47]), .B(IN_plaintext[47]), .S(IN_reset), .Z(
        LED_128_Instance_state1[47]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_48_U1 ( .A(
        LED_128_Instance_state0[48]), .B(IN_plaintext[48]), .S(IN_reset), .Z(
        LED_128_Instance_state1[48]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_49_U1 ( .A(
        LED_128_Instance_state0[49]), .B(IN_plaintext[49]), .S(IN_reset), .Z(
        LED_128_Instance_state1[49]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_50_U1 ( .A(
        LED_128_Instance_state0[50]), .B(IN_plaintext[50]), .S(IN_reset), .Z(
        LED_128_Instance_state1[50]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_51_U1 ( .A(
        LED_128_Instance_state0[51]), .B(IN_plaintext[51]), .S(IN_reset), .Z(
        LED_128_Instance_state1[51]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_52_U1 ( .A(
        LED_128_Instance_state0[52]), .B(IN_plaintext[52]), .S(IN_reset), .Z(
        LED_128_Instance_state1[52]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_53_U1 ( .A(
        LED_128_Instance_state0[53]), .B(IN_plaintext[53]), .S(IN_reset), .Z(
        LED_128_Instance_state1[53]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_54_U1 ( .A(
        LED_128_Instance_state0[54]), .B(IN_plaintext[54]), .S(IN_reset), .Z(
        LED_128_Instance_state1[54]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_55_U1 ( .A(
        LED_128_Instance_state0[55]), .B(IN_plaintext[55]), .S(IN_reset), .Z(
        LED_128_Instance_state1[55]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_56_U1 ( .A(
        LED_128_Instance_state0[56]), .B(IN_plaintext[56]), .S(IN_reset), .Z(
        LED_128_Instance_state1[56]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_57_U1 ( .A(
        LED_128_Instance_state0[57]), .B(IN_plaintext[57]), .S(IN_reset), .Z(
        LED_128_Instance_state1[57]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_58_U1 ( .A(
        LED_128_Instance_state0[58]), .B(IN_plaintext[58]), .S(IN_reset), .Z(
        LED_128_Instance_state1[58]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_59_U1 ( .A(
        LED_128_Instance_state0[59]), .B(IN_plaintext[59]), .S(IN_reset), .Z(
        LED_128_Instance_state1[59]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_60_U1 ( .A(
        LED_128_Instance_state0[60]), .B(IN_plaintext[60]), .S(IN_reset), .Z(
        LED_128_Instance_state1[60]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_61_U1 ( .A(
        LED_128_Instance_state0[61]), .B(IN_plaintext[61]), .S(IN_reset), .Z(
        LED_128_Instance_state1[61]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_62_U1 ( .A(
        LED_128_Instance_state0[62]), .B(IN_plaintext[62]), .S(IN_reset), .Z(
        LED_128_Instance_state1[62]) );
  MUX2_X1 LED_128_Instance_MUX_state1_mux_inst_63_U1 ( .A(
        LED_128_Instance_state0[63]), .B(IN_plaintext[63]), .S(IN_reset), .Z(
        LED_128_Instance_state1[63]) );
  INV_X1 LED_128_Instance_MUX_current_roundkey_U4 ( .A(
        LED_128_Instance_MUX_current_roundkey_n10), .ZN(
        LED_128_Instance_MUX_current_roundkey_n9) );
  INV_X1 LED_128_Instance_MUX_current_roundkey_U3 ( .A(LED_128_Instance_n12), 
        .ZN(LED_128_Instance_MUX_current_roundkey_n10) );
  INV_X1 LED_128_Instance_MUX_current_roundkey_U2 ( .A(
        LED_128_Instance_MUX_current_roundkey_n10), .ZN(
        LED_128_Instance_MUX_current_roundkey_n7) );
  INV_X1 LED_128_Instance_MUX_current_roundkey_U1 ( .A(
        LED_128_Instance_MUX_current_roundkey_n10), .ZN(
        LED_128_Instance_MUX_current_roundkey_n8) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1 ( .A(IN_key[64]), 
        .B(IN_key[0]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[0]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1 ( .A(IN_key[65]), 
        .B(IN_key[1]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[1]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1 ( .A(IN_key[66]), 
        .B(IN_key[2]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[2]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1 ( .A(IN_key[67]), 
        .B(IN_key[3]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[3]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1 ( .A(IN_key[68]), 
        .B(IN_key[4]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[4]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1 ( .A(IN_key[69]), 
        .B(IN_key[5]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[5]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1 ( .A(IN_key[70]), 
        .B(IN_key[6]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[6]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1 ( .A(IN_key[71]), 
        .B(IN_key[7]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[7]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1 ( .A(IN_key[72]), 
        .B(IN_key[8]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[8]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1 ( .A(IN_key[73]), 
        .B(IN_key[9]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[9]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1 ( .A(IN_key[74]), .B(IN_key[10]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[10]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1 ( .A(IN_key[75]), .B(IN_key[11]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[11]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1 ( .A(IN_key[76]), .B(IN_key[12]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[12]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1 ( .A(IN_key[77]), .B(IN_key[13]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[13]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1 ( .A(IN_key[78]), .B(IN_key[14]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[14]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1 ( .A(IN_key[79]), .B(IN_key[15]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[15]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1 ( .A(IN_key[80]), .B(IN_key[16]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[16]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1 ( .A(IN_key[81]), .B(IN_key[17]), .S(LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[17]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1 ( .A(IN_key[82]), .B(IN_key[18]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[18]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1 ( .A(IN_key[83]), .B(IN_key[19]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[19]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1 ( .A(IN_key[84]), .B(IN_key[20]), .S(LED_128_Instance_MUX_current_roundkey_n9), .Z(
        LED_128_Instance_current_roundkey[20]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1 ( .A(IN_key[85]), .B(IN_key[21]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[21]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1 ( .A(IN_key[86]), .B(IN_key[22]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[22]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1 ( .A(IN_key[87]), .B(IN_key[23]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[23]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1 ( .A(IN_key[88]), .B(IN_key[24]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[24]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1 ( .A(IN_key[89]), .B(IN_key[25]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[25]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1 ( .A(IN_key[90]), .B(IN_key[26]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[26]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1 ( .A(IN_key[91]), .B(IN_key[27]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[27]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1 ( .A(IN_key[92]), .B(IN_key[28]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[28]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1 ( .A(IN_key[93]), .B(IN_key[29]), .S(LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[29]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1 ( .A(IN_key[94]), .B(IN_key[30]), .S(LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[30]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1 ( .A(IN_key[95]), .B(IN_key[31]), .S(LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[31]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1 ( .A(IN_key[96]), .B(IN_key[32]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[32]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1 ( .A(IN_key[97]), .B(IN_key[33]), .S(LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[33]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1 ( .A(IN_key[98]), .B(IN_key[34]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[34]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1 ( .A(IN_key[99]), .B(IN_key[35]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[35]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1 ( .A(
        IN_key[100]), .B(IN_key[36]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[36]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1 ( .A(
        IN_key[101]), .B(IN_key[37]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[37]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1 ( .A(
        IN_key[102]), .B(IN_key[38]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[38]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1 ( .A(
        IN_key[103]), .B(IN_key[39]), .S(LED_128_Instance_n12), .Z(
        LED_128_Instance_current_roundkey[39]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1 ( .A(
        IN_key[104]), .B(IN_key[40]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[40]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1 ( .A(
        IN_key[105]), .B(IN_key[41]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[41]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1 ( .A(
        IN_key[106]), .B(IN_key[42]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[42]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1 ( .A(
        IN_key[107]), .B(IN_key[43]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[43]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1 ( .A(
        IN_key[108]), .B(IN_key[44]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[44]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1 ( .A(
        IN_key[109]), .B(IN_key[45]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[45]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1 ( .A(
        IN_key[110]), .B(IN_key[46]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[46]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1 ( .A(
        IN_key[111]), .B(IN_key[47]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[47]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1 ( .A(
        IN_key[112]), .B(IN_key[48]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[48]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1 ( .A(
        IN_key[113]), .B(IN_key[49]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[49]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1 ( .A(
        IN_key[114]), .B(IN_key[50]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[50]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1 ( .A(
        IN_key[115]), .B(IN_key[51]), .S(
        LED_128_Instance_MUX_current_roundkey_n8), .Z(
        LED_128_Instance_current_roundkey[51]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1 ( .A(
        IN_key[116]), .B(IN_key[52]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[52]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1 ( .A(
        IN_key[117]), .B(IN_key[53]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[53]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1 ( .A(
        IN_key[118]), .B(IN_key[54]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[54]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1 ( .A(
        IN_key[119]), .B(IN_key[55]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[55]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1 ( .A(
        IN_key[120]), .B(IN_key[56]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[56]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1 ( .A(
        IN_key[121]), .B(IN_key[57]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[57]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1 ( .A(
        IN_key[122]), .B(IN_key[58]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[58]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1 ( .A(
        IN_key[123]), .B(IN_key[59]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[59]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1 ( .A(
        IN_key[124]), .B(IN_key[60]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[60]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1 ( .A(
        IN_key[125]), .B(IN_key[61]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[61]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1 ( .A(
        IN_key[126]), .B(IN_key[62]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[62]) );
  MUX2_X1 LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1 ( .A(
        IN_key[127]), .B(IN_key[63]), .S(
        LED_128_Instance_MUX_current_roundkey_n7), .Z(
        LED_128_Instance_current_roundkey[63]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U64 ( .A(OUT_ciphertext[9]), 
        .B(LED_128_Instance_current_roundkey[9]), .Z(
        LED_128_Instance_addroundkey_tmp[9]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U63 ( .A(OUT_ciphertext[8]), 
        .B(LED_128_Instance_current_roundkey[8]), .Z(
        LED_128_Instance_addroundkey_tmp[8]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U62 ( .A(OUT_ciphertext[7]), 
        .B(LED_128_Instance_current_roundkey[7]), .Z(
        LED_128_Instance_addroundkey_tmp[7]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U61 ( .A(OUT_ciphertext[6]), 
        .B(LED_128_Instance_current_roundkey[6]), .Z(
        LED_128_Instance_addroundkey_tmp[6]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U60 ( .A(OUT_ciphertext[63]), 
        .B(LED_128_Instance_current_roundkey[63]), .Z(
        LED_128_Instance_addroundkey_tmp[63]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U59 ( .A(OUT_ciphertext[62]), 
        .B(LED_128_Instance_current_roundkey[62]), .Z(
        LED_128_Instance_addroundkey_tmp[62]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U58 ( .A(OUT_ciphertext[61]), 
        .B(LED_128_Instance_current_roundkey[61]), .Z(
        LED_128_Instance_addroundkey_tmp[61]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U57 ( .A(OUT_ciphertext[60]), 
        .B(LED_128_Instance_current_roundkey[60]), .Z(
        LED_128_Instance_addroundkey_tmp[60]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U56 ( .A(OUT_ciphertext[5]), 
        .B(LED_128_Instance_current_roundkey[5]), .Z(
        LED_128_Instance_addroundkey_tmp[5]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U55 ( .A(OUT_ciphertext[59]), 
        .B(LED_128_Instance_current_roundkey[59]), .Z(
        LED_128_Instance_addroundkey_tmp[59]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U54 ( .A(OUT_ciphertext[58]), 
        .B(LED_128_Instance_current_roundkey[58]), .Z(
        LED_128_Instance_addroundkey_tmp[58]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U53 ( .A(OUT_ciphertext[57]), 
        .B(LED_128_Instance_current_roundkey[57]), .Z(
        LED_128_Instance_addroundkey_tmp[57]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U52 ( .A(OUT_ciphertext[56]), 
        .B(LED_128_Instance_current_roundkey[56]), .Z(
        LED_128_Instance_addroundkey_tmp[56]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U51 ( .A(OUT_ciphertext[55]), 
        .B(LED_128_Instance_current_roundkey[55]), .Z(
        LED_128_Instance_addroundkey_tmp[55]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U50 ( .A(OUT_ciphertext[54]), 
        .B(LED_128_Instance_current_roundkey[54]), .Z(
        LED_128_Instance_addroundkey_tmp[54]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U49 ( .A(OUT_ciphertext[53]), 
        .B(LED_128_Instance_current_roundkey[53]), .Z(
        LED_128_Instance_addroundkey_tmp[53]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U48 ( .A(OUT_ciphertext[52]), 
        .B(LED_128_Instance_current_roundkey[52]), .Z(
        LED_128_Instance_addroundkey_tmp[52]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U47 ( .A(OUT_ciphertext[51]), 
        .B(LED_128_Instance_current_roundkey[51]), .Z(
        LED_128_Instance_addroundkey_tmp[51]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U46 ( .A(OUT_ciphertext[50]), 
        .B(LED_128_Instance_current_roundkey[50]), .Z(
        LED_128_Instance_addroundkey_tmp[50]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U45 ( .A(OUT_ciphertext[4]), 
        .B(LED_128_Instance_current_roundkey[4]), .Z(
        LED_128_Instance_addroundkey_tmp[4]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U44 ( .A(OUT_ciphertext[49]), 
        .B(LED_128_Instance_current_roundkey[49]), .Z(
        LED_128_Instance_addroundkey_tmp[49]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U43 ( .A(OUT_ciphertext[48]), 
        .B(LED_128_Instance_current_roundkey[48]), .Z(
        LED_128_Instance_addroundkey_tmp[48]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U42 ( .A(OUT_ciphertext[47]), 
        .B(LED_128_Instance_current_roundkey[47]), .Z(
        LED_128_Instance_addroundkey_tmp[47]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U41 ( .A(OUT_ciphertext[46]), 
        .B(LED_128_Instance_current_roundkey[46]), .Z(
        LED_128_Instance_addroundkey_tmp[46]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U40 ( .A(OUT_ciphertext[45]), 
        .B(LED_128_Instance_current_roundkey[45]), .Z(
        LED_128_Instance_addroundkey_tmp[45]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U39 ( .A(OUT_ciphertext[44]), 
        .B(LED_128_Instance_current_roundkey[44]), .Z(
        LED_128_Instance_addroundkey_tmp[44]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U38 ( .A(OUT_ciphertext[43]), 
        .B(LED_128_Instance_current_roundkey[43]), .Z(
        LED_128_Instance_addroundkey_tmp[43]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U37 ( .A(OUT_ciphertext[42]), 
        .B(LED_128_Instance_current_roundkey[42]), .Z(
        LED_128_Instance_addroundkey_tmp[42]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U36 ( .A(OUT_ciphertext[41]), 
        .B(LED_128_Instance_current_roundkey[41]), .Z(
        LED_128_Instance_addroundkey_tmp[41]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U35 ( .A(OUT_ciphertext[40]), 
        .B(LED_128_Instance_current_roundkey[40]), .Z(
        LED_128_Instance_addroundkey_tmp[40]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U34 ( .A(OUT_ciphertext[3]), 
        .B(LED_128_Instance_current_roundkey[3]), .Z(
        LED_128_Instance_addroundkey_tmp[3]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U33 ( .A(OUT_ciphertext[39]), 
        .B(LED_128_Instance_current_roundkey[39]), .Z(
        LED_128_Instance_addroundkey_tmp[39]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U32 ( .A(OUT_ciphertext[38]), 
        .B(LED_128_Instance_current_roundkey[38]), .Z(
        LED_128_Instance_addroundkey_tmp[38]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U31 ( .A(OUT_ciphertext[37]), 
        .B(LED_128_Instance_current_roundkey[37]), .Z(
        LED_128_Instance_addroundkey_tmp[37]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U30 ( .A(OUT_ciphertext[36]), 
        .B(LED_128_Instance_current_roundkey[36]), .Z(
        LED_128_Instance_addroundkey_tmp[36]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U29 ( .A(OUT_ciphertext[35]), 
        .B(LED_128_Instance_current_roundkey[35]), .Z(
        LED_128_Instance_addroundkey_tmp[35]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U28 ( .A(OUT_ciphertext[34]), 
        .B(LED_128_Instance_current_roundkey[34]), .Z(
        LED_128_Instance_addroundkey_tmp[34]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U27 ( .A(OUT_ciphertext[33]), 
        .B(LED_128_Instance_current_roundkey[33]), .Z(
        LED_128_Instance_addroundkey_tmp[33]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U26 ( .A(OUT_ciphertext[32]), 
        .B(LED_128_Instance_current_roundkey[32]), .Z(
        LED_128_Instance_addroundkey_tmp[32]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U25 ( .A(OUT_ciphertext[31]), 
        .B(LED_128_Instance_current_roundkey[31]), .Z(
        LED_128_Instance_addroundkey_tmp[31]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U24 ( .A(OUT_ciphertext[30]), 
        .B(LED_128_Instance_current_roundkey[30]), .Z(
        LED_128_Instance_addroundkey_tmp[30]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U23 ( .A(OUT_ciphertext[2]), 
        .B(LED_128_Instance_current_roundkey[2]), .Z(
        LED_128_Instance_addroundkey_tmp[2]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U22 ( .A(OUT_ciphertext[29]), 
        .B(LED_128_Instance_current_roundkey[29]), .Z(
        LED_128_Instance_addroundkey_tmp[29]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U21 ( .A(OUT_ciphertext[28]), 
        .B(LED_128_Instance_current_roundkey[28]), .Z(
        LED_128_Instance_addroundkey_tmp[28]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U20 ( .A(OUT_ciphertext[27]), 
        .B(LED_128_Instance_current_roundkey[27]), .Z(
        LED_128_Instance_addroundkey_tmp[27]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U19 ( .A(OUT_ciphertext[26]), 
        .B(LED_128_Instance_current_roundkey[26]), .Z(
        LED_128_Instance_addroundkey_tmp[26]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U18 ( .A(OUT_ciphertext[25]), 
        .B(LED_128_Instance_current_roundkey[25]), .Z(
        LED_128_Instance_addroundkey_tmp[25]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U17 ( .A(OUT_ciphertext[24]), 
        .B(LED_128_Instance_current_roundkey[24]), .Z(
        LED_128_Instance_addroundkey_tmp[24]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U16 ( .A(OUT_ciphertext[23]), 
        .B(LED_128_Instance_current_roundkey[23]), .Z(
        LED_128_Instance_addroundkey_tmp[23]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U15 ( .A(OUT_ciphertext[22]), 
        .B(LED_128_Instance_current_roundkey[22]), .Z(
        LED_128_Instance_addroundkey_tmp[22]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U14 ( .A(OUT_ciphertext[21]), 
        .B(LED_128_Instance_current_roundkey[21]), .Z(
        LED_128_Instance_addroundkey_tmp[21]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U13 ( .A(OUT_ciphertext[20]), 
        .B(LED_128_Instance_current_roundkey[20]), .Z(
        LED_128_Instance_addroundkey_tmp[20]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U12 ( .A(OUT_ciphertext[1]), 
        .B(LED_128_Instance_current_roundkey[1]), .Z(
        LED_128_Instance_addroundkey_tmp[1]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U11 ( .A(OUT_ciphertext[19]), 
        .B(LED_128_Instance_current_roundkey[19]), .Z(
        LED_128_Instance_addroundkey_tmp[19]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U10 ( .A(OUT_ciphertext[18]), 
        .B(LED_128_Instance_current_roundkey[18]), .Z(
        LED_128_Instance_addroundkey_tmp[18]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U9 ( .A(OUT_ciphertext[17]), 
        .B(LED_128_Instance_current_roundkey[17]), .Z(
        LED_128_Instance_addroundkey_tmp[17]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U8 ( .A(OUT_ciphertext[16]), 
        .B(LED_128_Instance_current_roundkey[16]), .Z(
        LED_128_Instance_addroundkey_tmp[16]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U7 ( .A(OUT_ciphertext[15]), 
        .B(LED_128_Instance_current_roundkey[15]), .Z(
        LED_128_Instance_addroundkey_tmp[15]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U6 ( .A(OUT_ciphertext[14]), 
        .B(LED_128_Instance_current_roundkey[14]), .Z(
        LED_128_Instance_addroundkey_tmp[14]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U5 ( .A(OUT_ciphertext[13]), 
        .B(LED_128_Instance_current_roundkey[13]), .Z(
        LED_128_Instance_addroundkey_tmp[13]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U4 ( .A(OUT_ciphertext[12]), 
        .B(LED_128_Instance_current_roundkey[12]), .Z(
        LED_128_Instance_addroundkey_tmp[12]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U3 ( .A(OUT_ciphertext[11]), 
        .B(LED_128_Instance_current_roundkey[11]), .Z(
        LED_128_Instance_addroundkey_tmp[11]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U2 ( .A(OUT_ciphertext[10]), 
        .B(LED_128_Instance_current_roundkey[10]), .Z(
        LED_128_Instance_addroundkey_tmp[10]) );
  XOR2_X1 LED_128_Instance_addRoundKey_instance_U1 ( .A(OUT_ciphertext[0]), 
        .B(LED_128_Instance_current_roundkey[0]), .Z(
        LED_128_Instance_addroundkey_tmp[0]) );
  INV_X2 LED_128_Instance_MUX_addroundkey_out_U3 ( .A(
        LED_128_Instance_MUX_addroundkey_out_n9), .ZN(
        LED_128_Instance_MUX_addroundkey_out_n7) );
  INV_X1 LED_128_Instance_MUX_addroundkey_out_U2 ( .A(LED_128_Instance_n31), 
        .ZN(LED_128_Instance_MUX_addroundkey_out_n9) );
  INV_X1 LED_128_Instance_MUX_addroundkey_out_U1 ( .A(
        LED_128_Instance_MUX_addroundkey_out_n9), .ZN(
        LED_128_Instance_MUX_addroundkey_out_n8) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1 ( .A(
        OUT_ciphertext[0]), .B(LED_128_Instance_addroundkey_tmp[0]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_0_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1 ( .A(
        OUT_ciphertext[1]), .B(LED_128_Instance_addroundkey_tmp[1]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_1_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1 ( .A(
        OUT_ciphertext[2]), .B(LED_128_Instance_addroundkey_tmp[2]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_2_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1 ( .A(
        OUT_ciphertext[3]), .B(LED_128_Instance_addroundkey_tmp[3]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_3_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1 ( .A(
        OUT_ciphertext[4]), .B(LED_128_Instance_addroundkey_tmp[4]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addroundkey_out_4_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1 ( .A(
        OUT_ciphertext[5]), .B(LED_128_Instance_addroundkey_tmp[5]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addroundkey_out_5_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1 ( .A(
        OUT_ciphertext[6]), .B(LED_128_Instance_addroundkey_tmp[6]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addroundkey_out_6_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1 ( .A(
        OUT_ciphertext[7]), .B(LED_128_Instance_addroundkey_tmp[7]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[7]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1 ( .A(
        OUT_ciphertext[8]), .B(LED_128_Instance_addroundkey_tmp[8]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[8]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1 ( .A(
        OUT_ciphertext[9]), .B(LED_128_Instance_addroundkey_tmp[9]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[9]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1 ( .A(
        OUT_ciphertext[10]), .B(LED_128_Instance_addroundkey_tmp[10]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[10]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1 ( .A(
        OUT_ciphertext[11]), .B(LED_128_Instance_addroundkey_tmp[11]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[11]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1 ( .A(
        OUT_ciphertext[12]), .B(LED_128_Instance_addroundkey_tmp[12]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[12]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1 ( .A(
        OUT_ciphertext[13]), .B(LED_128_Instance_addroundkey_tmp[13]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[13]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1 ( .A(
        OUT_ciphertext[14]), .B(LED_128_Instance_addroundkey_tmp[14]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[14]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1 ( .A(
        OUT_ciphertext[15]), .B(LED_128_Instance_addroundkey_tmp[15]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addconst_out[15]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1 ( .A(
        OUT_ciphertext[16]), .B(LED_128_Instance_addroundkey_tmp[16]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_16_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1 ( .A(
        OUT_ciphertext[17]), .B(LED_128_Instance_addroundkey_tmp[17]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_17_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1 ( .A(
        OUT_ciphertext[18]), .B(LED_128_Instance_addroundkey_tmp[18]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_18_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1 ( .A(
        OUT_ciphertext[19]), .B(LED_128_Instance_addroundkey_tmp[19]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_19_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1 ( .A(
        OUT_ciphertext[20]), .B(LED_128_Instance_addroundkey_tmp[20]), .S(
        LED_128_Instance_MUX_addroundkey_out_n8), .Z(
        LED_128_Instance_addroundkey_out_20_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1 ( .A(
        OUT_ciphertext[21]), .B(LED_128_Instance_addroundkey_tmp[21]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_21_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1 ( .A(
        OUT_ciphertext[22]), .B(LED_128_Instance_addroundkey_tmp[22]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_22_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1 ( .A(
        OUT_ciphertext[23]), .B(LED_128_Instance_addroundkey_tmp[23]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addconst_out[23]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1 ( .A(
        OUT_ciphertext[24]), .B(LED_128_Instance_addroundkey_tmp[24]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addconst_out[24]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1 ( .A(
        OUT_ciphertext[25]), .B(LED_128_Instance_addroundkey_tmp[25]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addconst_out[25]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1 ( .A(
        OUT_ciphertext[26]), .B(LED_128_Instance_addroundkey_tmp[26]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addconst_out[26]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1 ( .A(
        OUT_ciphertext[27]), .B(LED_128_Instance_addroundkey_tmp[27]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addconst_out[27]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1 ( .A(
        OUT_ciphertext[28]), .B(LED_128_Instance_addroundkey_tmp[28]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[28]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1 ( .A(
        OUT_ciphertext[29]), .B(LED_128_Instance_addroundkey_tmp[29]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[29]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1 ( .A(
        OUT_ciphertext[30]), .B(LED_128_Instance_addroundkey_tmp[30]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[30]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1 ( .A(
        OUT_ciphertext[31]), .B(LED_128_Instance_addroundkey_tmp[31]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[31]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1 ( .A(
        OUT_ciphertext[32]), .B(LED_128_Instance_addroundkey_tmp[32]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_32_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1 ( .A(
        OUT_ciphertext[33]), .B(LED_128_Instance_addroundkey_tmp[33]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_33_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1 ( .A(
        OUT_ciphertext[34]), .B(LED_128_Instance_addroundkey_tmp[34]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_34_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1 ( .A(
        OUT_ciphertext[35]), .B(LED_128_Instance_addroundkey_tmp[35]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_35_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1 ( .A(
        OUT_ciphertext[36]), .B(LED_128_Instance_addroundkey_tmp[36]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_36_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1 ( .A(
        OUT_ciphertext[37]), .B(LED_128_Instance_addroundkey_tmp[37]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_37_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1 ( .A(
        OUT_ciphertext[38]), .B(LED_128_Instance_addroundkey_tmp[38]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_38_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1 ( .A(
        OUT_ciphertext[39]), .B(LED_128_Instance_addroundkey_tmp[39]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[39]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1 ( .A(
        OUT_ciphertext[40]), .B(LED_128_Instance_addroundkey_tmp[40]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[40]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1 ( .A(
        OUT_ciphertext[41]), .B(LED_128_Instance_addroundkey_tmp[41]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[41]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1 ( .A(
        OUT_ciphertext[42]), .B(LED_128_Instance_addroundkey_tmp[42]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[42]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1 ( .A(
        OUT_ciphertext[43]), .B(LED_128_Instance_addroundkey_tmp[43]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[43]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1 ( .A(
        OUT_ciphertext[44]), .B(LED_128_Instance_addroundkey_tmp[44]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[44]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1 ( .A(
        OUT_ciphertext[45]), .B(LED_128_Instance_addroundkey_tmp[45]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[45]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1 ( .A(
        OUT_ciphertext[46]), .B(LED_128_Instance_addroundkey_tmp[46]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[46]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1 ( .A(
        OUT_ciphertext[47]), .B(LED_128_Instance_addroundkey_tmp[47]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[47]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1 ( .A(
        OUT_ciphertext[48]), .B(LED_128_Instance_addroundkey_tmp[48]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_48_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1 ( .A(
        OUT_ciphertext[49]), .B(LED_128_Instance_addroundkey_tmp[49]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_49_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1 ( .A(
        OUT_ciphertext[50]), .B(LED_128_Instance_addroundkey_tmp[50]), .S(
        LED_128_Instance_n31), .Z(LED_128_Instance_addroundkey_out_50_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1 ( .A(
        OUT_ciphertext[51]), .B(LED_128_Instance_addroundkey_tmp[51]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_51_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1 ( .A(
        OUT_ciphertext[52]), .B(LED_128_Instance_addroundkey_tmp[52]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_52_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1 ( .A(
        OUT_ciphertext[53]), .B(LED_128_Instance_addroundkey_tmp[53]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_53_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1 ( .A(
        OUT_ciphertext[54]), .B(LED_128_Instance_addroundkey_tmp[54]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addroundkey_out_54_) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1 ( .A(
        OUT_ciphertext[55]), .B(LED_128_Instance_addroundkey_tmp[55]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[55]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1 ( .A(
        OUT_ciphertext[56]), .B(LED_128_Instance_addroundkey_tmp[56]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[56]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1 ( .A(
        OUT_ciphertext[57]), .B(LED_128_Instance_addroundkey_tmp[57]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[57]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1 ( .A(
        OUT_ciphertext[58]), .B(LED_128_Instance_addroundkey_tmp[58]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[58]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1 ( .A(
        OUT_ciphertext[59]), .B(LED_128_Instance_addroundkey_tmp[59]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[59]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1 ( .A(
        OUT_ciphertext[60]), .B(LED_128_Instance_addroundkey_tmp[60]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[60]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1 ( .A(
        OUT_ciphertext[61]), .B(LED_128_Instance_addroundkey_tmp[61]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[61]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1 ( .A(
        OUT_ciphertext[62]), .B(LED_128_Instance_addroundkey_tmp[62]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[62]) );
  MUX2_X1 LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1 ( .A(
        OUT_ciphertext[63]), .B(LED_128_Instance_addroundkey_tmp[63]), .S(
        LED_128_Instance_MUX_addroundkey_out_n7), .Z(
        LED_128_Instance_addconst_out[63]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U28 ( .A(roundconstant[5]), 
        .B(LED_128_Instance_addroundkey_out_6_), .Z(
        LED_128_Instance_addconst_out[6]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U27 ( .A(roundconstant[4]), 
        .B(LED_128_Instance_addroundkey_out_5_), .Z(
        LED_128_Instance_addconst_out[5]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U26 ( .A(roundconstant[2]), 
        .B(LED_128_Instance_addroundkey_out_54_), .Z(
        LED_128_Instance_addconst_out[54]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U25 ( .A(roundconstant[1]), 
        .B(LED_128_Instance_addroundkey_out_53_), .Z(
        LED_128_Instance_addconst_out[53]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U24 ( .A(roundconstant[0]), 
        .B(LED_128_Instance_addroundkey_out_52_), .Z(
        LED_128_Instance_addconst_out[52]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U23 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_51_), .Z(
        LED_128_Instance_addconst_out[51]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U22 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_50_), .Z(
        LED_128_Instance_addconst_out[50]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U21 ( .A(roundconstant[3]), 
        .B(LED_128_Instance_addroundkey_out_4_), .Z(
        LED_128_Instance_addconst_out[4]) );
  XNOR2_X1 LED_128_Instance_AddConstants_instance_U20 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_49_), .ZN(
        LED_128_Instance_addconst_out[49]) );
  XNOR2_X1 LED_128_Instance_AddConstants_instance_U19 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_48_), .ZN(
        LED_128_Instance_addconst_out[48]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U18 ( .A(1'b1), .B(
        LED_128_Instance_addroundkey_out_3_), .Z(
        LED_128_Instance_addconst_out[3]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U17 ( .A(roundconstant[5]), 
        .B(LED_128_Instance_addroundkey_out_38_), .Z(
        LED_128_Instance_addconst_out[38]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U16 ( .A(roundconstant[4]), 
        .B(LED_128_Instance_addroundkey_out_37_), .Z(
        LED_128_Instance_addconst_out[37]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U15 ( .A(roundconstant[3]), 
        .B(LED_128_Instance_addroundkey_out_36_), .Z(
        LED_128_Instance_addconst_out[36]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U14 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_35_), .Z(
        LED_128_Instance_addconst_out[35]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U13 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_34_), .Z(
        LED_128_Instance_addconst_out[34]) );
  XNOR2_X1 LED_128_Instance_AddConstants_instance_U12 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_33_), .ZN(
        LED_128_Instance_addconst_out[33]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U11 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_32_), .Z(
        LED_128_Instance_addconst_out[32]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U10 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_2_), .Z(
        LED_128_Instance_addconst_out[2]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U9 ( .A(roundconstant[2]), 
        .B(LED_128_Instance_addroundkey_out_22_), .Z(
        LED_128_Instance_addconst_out[22]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U8 ( .A(roundconstant[1]), 
        .B(LED_128_Instance_addroundkey_out_21_), .Z(
        LED_128_Instance_addconst_out[21]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U7 ( .A(roundconstant[0]), 
        .B(LED_128_Instance_addroundkey_out_20_), .Z(
        LED_128_Instance_addconst_out[20]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U6 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_1_), .Z(
        LED_128_Instance_addconst_out[1]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U5 ( .A(1'b1), .B(
        LED_128_Instance_addroundkey_out_19_), .Z(
        LED_128_Instance_addconst_out[19]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U4 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_18_), .Z(
        LED_128_Instance_addconst_out[18]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U3 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_17_), .Z(
        LED_128_Instance_addconst_out[17]) );
  XNOR2_X1 LED_128_Instance_AddConstants_instance_U2 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_16_), .ZN(
        LED_128_Instance_addconst_out[16]) );
  XOR2_X1 LED_128_Instance_AddConstants_instance_U1 ( .A(1'b0), .B(
        LED_128_Instance_addroundkey_out_0_), .Z(
        LED_128_Instance_addconst_out[0]) );
  INV_X1 LED_128_Instance_SBox_Instance_0_U3 ( .A(
        LED_128_Instance_SBox_Instance_0_L0), .ZN(
        LED_128_Instance_SBox_Instance_0_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_0_U2 ( .A(
        LED_128_Instance_addconst_out[3]), .ZN(
        LED_128_Instance_SBox_Instance_0_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_0_U1 ( .A(
        LED_128_Instance_addconst_out[1]), .ZN(
        LED_128_Instance_SBox_Instance_0_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[2]), .B(LED_128_Instance_addconst_out[1]), .Z(LED_128_Instance_SBox_Instance_0_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[1]), .B(LED_128_Instance_addconst_out[0]), .Z(LED_128_Instance_SBox_Instance_0_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L1), .B(
        LED_128_Instance_addconst_out[3]), .Z(
        LED_128_Instance_SBox_Instance_0_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_T0), .B(
        LED_128_Instance_SBox_Instance_0_L2), .ZN(
        LED_128_Instance_SBox_Instance_0_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[3]), .B(LED_128_Instance_addconst_out[0]), .Z(LED_128_Instance_SBox_Instance_0_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L3), .B(
        LED_128_Instance_SBox_Instance_0_L0), .Z(
        LED_128_Instance_SBox_Instance_0_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[3]), .B(LED_128_Instance_addconst_out[1]), .Z(LED_128_Instance_SBox_Instance_0_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_T0), .B(
        LED_128_Instance_SBox_Instance_0_T2), .Z(
        LED_128_Instance_SBox_Instance_0_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L4), .B(
        LED_128_Instance_SBox_Instance_0_L5), .ZN(
        LED_128_Instance_SBox_Instance_0_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L1), .B(
        LED_128_Instance_addconst_out[2]), .Z(
        LED_128_Instance_SBox_Instance_0_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_0_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_0_n1), .A2(
        LED_128_Instance_SBox_Instance_0_n2), .ZN(
        LED_128_Instance_SBox_Instance_0_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_0_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_0_Q2), .A2(
        LED_128_Instance_SBox_Instance_0_Q3), .ZN(
        LED_128_Instance_SBox_Instance_0_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_0_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_0_n3), .A2(
        LED_128_Instance_addconst_out[2]), .ZN(
        LED_128_Instance_SBox_Instance_0_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_0_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_0_Q6), .A2(
        LED_128_Instance_SBox_Instance_0_Q7), .ZN(
        LED_128_Instance_SBox_Instance_0_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L5), .B(
        LED_128_Instance_SBox_Instance_0_T3), .Z(
        LED_128_Instance_SBox_Instance_0_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[0]), .B(
        LED_128_Instance_SBox_Instance_0_L7), .Z(
        LED_128_Instance_subcells_out[3]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L5), .B(
        LED_128_Instance_SBox_Instance_0_T1), .Z(
        LED_128_Instance_SBox_Instance_0_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L1), .B(
        LED_128_Instance_SBox_Instance_0_L8), .Z(
        LED_128_Instance_subcells_out[2]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L4), .B(
        LED_128_Instance_SBox_Instance_0_T3), .Z(
        LED_128_Instance_subcells_out[1]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_0_L3), .B(
        LED_128_Instance_SBox_Instance_0_T2), .Z(
        LED_128_Instance_subcells_out[0]) );
  INV_X1 LED_128_Instance_SBox_Instance_1_U3 ( .A(
        LED_128_Instance_SBox_Instance_1_L0), .ZN(
        LED_128_Instance_SBox_Instance_1_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_1_U2 ( .A(
        LED_128_Instance_addconst_out[7]), .ZN(
        LED_128_Instance_SBox_Instance_1_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_1_U1 ( .A(
        LED_128_Instance_addconst_out[5]), .ZN(
        LED_128_Instance_SBox_Instance_1_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[6]), .B(LED_128_Instance_addconst_out[5]), .Z(LED_128_Instance_SBox_Instance_1_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[5]), .B(LED_128_Instance_addconst_out[4]), .Z(LED_128_Instance_SBox_Instance_1_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L1), .B(
        LED_128_Instance_addconst_out[7]), .Z(
        LED_128_Instance_SBox_Instance_1_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_T0), .B(
        LED_128_Instance_SBox_Instance_1_L2), .ZN(
        LED_128_Instance_SBox_Instance_1_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[7]), .B(LED_128_Instance_addconst_out[4]), .Z(LED_128_Instance_SBox_Instance_1_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L3), .B(
        LED_128_Instance_SBox_Instance_1_L0), .Z(
        LED_128_Instance_SBox_Instance_1_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[7]), .B(LED_128_Instance_addconst_out[5]), .Z(LED_128_Instance_SBox_Instance_1_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_T0), .B(
        LED_128_Instance_SBox_Instance_1_T2), .Z(
        LED_128_Instance_SBox_Instance_1_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L4), .B(
        LED_128_Instance_SBox_Instance_1_L5), .ZN(
        LED_128_Instance_SBox_Instance_1_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L1), .B(
        LED_128_Instance_addconst_out[6]), .Z(
        LED_128_Instance_SBox_Instance_1_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_1_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_1_n1), .A2(
        LED_128_Instance_SBox_Instance_1_n2), .ZN(
        LED_128_Instance_SBox_Instance_1_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_1_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_1_Q2), .A2(
        LED_128_Instance_SBox_Instance_1_Q3), .ZN(
        LED_128_Instance_SBox_Instance_1_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_1_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_1_n3), .A2(
        LED_128_Instance_addconst_out[6]), .ZN(
        LED_128_Instance_SBox_Instance_1_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_1_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_1_Q6), .A2(
        LED_128_Instance_SBox_Instance_1_Q7), .ZN(
        LED_128_Instance_SBox_Instance_1_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L5), .B(
        LED_128_Instance_SBox_Instance_1_T3), .Z(
        LED_128_Instance_SBox_Instance_1_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[4]), .B(
        LED_128_Instance_SBox_Instance_1_L7), .Z(
        LED_128_Instance_subcells_out[7]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L5), .B(
        LED_128_Instance_SBox_Instance_1_T1), .Z(
        LED_128_Instance_SBox_Instance_1_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L1), .B(
        LED_128_Instance_SBox_Instance_1_L8), .Z(
        LED_128_Instance_subcells_out[6]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L4), .B(
        LED_128_Instance_SBox_Instance_1_T3), .Z(
        LED_128_Instance_subcells_out[5]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_1_L3), .B(
        LED_128_Instance_SBox_Instance_1_T2), .Z(
        LED_128_Instance_subcells_out[4]) );
  INV_X1 LED_128_Instance_SBox_Instance_2_U3 ( .A(
        LED_128_Instance_SBox_Instance_2_L0), .ZN(
        LED_128_Instance_SBox_Instance_2_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_2_U2 ( .A(
        LED_128_Instance_addconst_out[11]), .ZN(
        LED_128_Instance_SBox_Instance_2_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_2_U1 ( .A(
        LED_128_Instance_addconst_out[9]), .ZN(
        LED_128_Instance_SBox_Instance_2_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[10]), .B(
        LED_128_Instance_addconst_out[9]), .Z(
        LED_128_Instance_SBox_Instance_2_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[9]), .B(LED_128_Instance_addconst_out[8]), .Z(LED_128_Instance_SBox_Instance_2_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L1), .B(
        LED_128_Instance_addconst_out[11]), .Z(
        LED_128_Instance_SBox_Instance_2_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_T0), .B(
        LED_128_Instance_SBox_Instance_2_L2), .ZN(
        LED_128_Instance_SBox_Instance_2_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[11]), .B(
        LED_128_Instance_addconst_out[8]), .Z(
        LED_128_Instance_SBox_Instance_2_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L3), .B(
        LED_128_Instance_SBox_Instance_2_L0), .Z(
        LED_128_Instance_SBox_Instance_2_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[11]), .B(
        LED_128_Instance_addconst_out[9]), .Z(
        LED_128_Instance_SBox_Instance_2_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_T0), .B(
        LED_128_Instance_SBox_Instance_2_T2), .Z(
        LED_128_Instance_SBox_Instance_2_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L4), .B(
        LED_128_Instance_SBox_Instance_2_L5), .ZN(
        LED_128_Instance_SBox_Instance_2_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L1), .B(
        LED_128_Instance_addconst_out[10]), .Z(
        LED_128_Instance_SBox_Instance_2_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_2_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_2_n1), .A2(
        LED_128_Instance_SBox_Instance_2_n2), .ZN(
        LED_128_Instance_SBox_Instance_2_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_2_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_2_Q2), .A2(
        LED_128_Instance_SBox_Instance_2_Q3), .ZN(
        LED_128_Instance_SBox_Instance_2_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_2_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_2_n3), .A2(
        LED_128_Instance_addconst_out[10]), .ZN(
        LED_128_Instance_SBox_Instance_2_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_2_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_2_Q6), .A2(
        LED_128_Instance_SBox_Instance_2_Q7), .ZN(
        LED_128_Instance_SBox_Instance_2_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L5), .B(
        LED_128_Instance_SBox_Instance_2_T3), .Z(
        LED_128_Instance_SBox_Instance_2_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[8]), .B(
        LED_128_Instance_SBox_Instance_2_L7), .Z(
        LED_128_Instance_subcells_out[11]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L5), .B(
        LED_128_Instance_SBox_Instance_2_T1), .Z(
        LED_128_Instance_SBox_Instance_2_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L1), .B(
        LED_128_Instance_SBox_Instance_2_L8), .Z(
        LED_128_Instance_subcells_out[10]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L4), .B(
        LED_128_Instance_SBox_Instance_2_T3), .Z(
        LED_128_Instance_subcells_out[9]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_2_L3), .B(
        LED_128_Instance_SBox_Instance_2_T2), .Z(
        LED_128_Instance_subcells_out[8]) );
  INV_X1 LED_128_Instance_SBox_Instance_3_U3 ( .A(
        LED_128_Instance_SBox_Instance_3_L0), .ZN(
        LED_128_Instance_SBox_Instance_3_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_3_U2 ( .A(
        LED_128_Instance_addconst_out[15]), .ZN(
        LED_128_Instance_SBox_Instance_3_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_3_U1 ( .A(
        LED_128_Instance_addconst_out[13]), .ZN(
        LED_128_Instance_SBox_Instance_3_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[14]), .B(
        LED_128_Instance_addconst_out[13]), .Z(
        LED_128_Instance_SBox_Instance_3_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[13]), .B(
        LED_128_Instance_addconst_out[12]), .Z(
        LED_128_Instance_SBox_Instance_3_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L1), .B(
        LED_128_Instance_addconst_out[15]), .Z(
        LED_128_Instance_SBox_Instance_3_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_T0), .B(
        LED_128_Instance_SBox_Instance_3_L2), .ZN(
        LED_128_Instance_SBox_Instance_3_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[15]), .B(
        LED_128_Instance_addconst_out[12]), .Z(
        LED_128_Instance_SBox_Instance_3_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L3), .B(
        LED_128_Instance_SBox_Instance_3_L0), .Z(
        LED_128_Instance_SBox_Instance_3_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[15]), .B(
        LED_128_Instance_addconst_out[13]), .Z(
        LED_128_Instance_SBox_Instance_3_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_T0), .B(
        LED_128_Instance_SBox_Instance_3_T2), .Z(
        LED_128_Instance_SBox_Instance_3_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L4), .B(
        LED_128_Instance_SBox_Instance_3_L5), .ZN(
        LED_128_Instance_SBox_Instance_3_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L1), .B(
        LED_128_Instance_addconst_out[14]), .Z(
        LED_128_Instance_SBox_Instance_3_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_3_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_3_n1), .A2(
        LED_128_Instance_SBox_Instance_3_n2), .ZN(
        LED_128_Instance_SBox_Instance_3_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_3_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_3_Q2), .A2(
        LED_128_Instance_SBox_Instance_3_Q3), .ZN(
        LED_128_Instance_SBox_Instance_3_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_3_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_3_n3), .A2(
        LED_128_Instance_addconst_out[14]), .ZN(
        LED_128_Instance_SBox_Instance_3_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_3_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_3_Q6), .A2(
        LED_128_Instance_SBox_Instance_3_Q7), .ZN(
        LED_128_Instance_SBox_Instance_3_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L5), .B(
        LED_128_Instance_SBox_Instance_3_T3), .Z(
        LED_128_Instance_SBox_Instance_3_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[12]), .B(
        LED_128_Instance_SBox_Instance_3_L7), .Z(
        LED_128_Instance_subcells_out[15]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L5), .B(
        LED_128_Instance_SBox_Instance_3_T1), .Z(
        LED_128_Instance_SBox_Instance_3_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L1), .B(
        LED_128_Instance_SBox_Instance_3_L8), .Z(
        LED_128_Instance_subcells_out[14]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L4), .B(
        LED_128_Instance_SBox_Instance_3_T3), .Z(
        LED_128_Instance_subcells_out[13]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_3_L3), .B(
        LED_128_Instance_SBox_Instance_3_T2), .Z(
        LED_128_Instance_subcells_out[12]) );
  INV_X1 LED_128_Instance_SBox_Instance_4_U3 ( .A(
        LED_128_Instance_SBox_Instance_4_L0), .ZN(
        LED_128_Instance_SBox_Instance_4_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_4_U2 ( .A(
        LED_128_Instance_addconst_out[19]), .ZN(
        LED_128_Instance_SBox_Instance_4_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_4_U1 ( .A(
        LED_128_Instance_addconst_out[17]), .ZN(
        LED_128_Instance_SBox_Instance_4_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[18]), .B(
        LED_128_Instance_addconst_out[17]), .Z(
        LED_128_Instance_SBox_Instance_4_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[17]), .B(
        LED_128_Instance_addconst_out[16]), .Z(
        LED_128_Instance_SBox_Instance_4_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L1), .B(
        LED_128_Instance_addconst_out[19]), .Z(
        LED_128_Instance_SBox_Instance_4_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_T0), .B(
        LED_128_Instance_SBox_Instance_4_L2), .ZN(
        LED_128_Instance_SBox_Instance_4_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[19]), .B(
        LED_128_Instance_addconst_out[16]), .Z(
        LED_128_Instance_SBox_Instance_4_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L3), .B(
        LED_128_Instance_SBox_Instance_4_L0), .Z(
        LED_128_Instance_SBox_Instance_4_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[19]), .B(
        LED_128_Instance_addconst_out[17]), .Z(
        LED_128_Instance_SBox_Instance_4_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_T0), .B(
        LED_128_Instance_SBox_Instance_4_T2), .Z(
        LED_128_Instance_SBox_Instance_4_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L4), .B(
        LED_128_Instance_SBox_Instance_4_L5), .ZN(
        LED_128_Instance_SBox_Instance_4_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L1), .B(
        LED_128_Instance_addconst_out[18]), .Z(
        LED_128_Instance_SBox_Instance_4_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_4_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_4_n1), .A2(
        LED_128_Instance_SBox_Instance_4_n2), .ZN(
        LED_128_Instance_SBox_Instance_4_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_4_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_4_Q2), .A2(
        LED_128_Instance_SBox_Instance_4_Q3), .ZN(
        LED_128_Instance_SBox_Instance_4_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_4_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_4_n3), .A2(
        LED_128_Instance_addconst_out[18]), .ZN(
        LED_128_Instance_SBox_Instance_4_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_4_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_4_Q6), .A2(
        LED_128_Instance_SBox_Instance_4_Q7), .ZN(
        LED_128_Instance_SBox_Instance_4_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L5), .B(
        LED_128_Instance_SBox_Instance_4_T3), .Z(
        LED_128_Instance_SBox_Instance_4_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[16]), .B(
        LED_128_Instance_SBox_Instance_4_L7), .Z(
        LED_128_Instance_subcells_out[19]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L5), .B(
        LED_128_Instance_SBox_Instance_4_T1), .Z(
        LED_128_Instance_SBox_Instance_4_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L1), .B(
        LED_128_Instance_SBox_Instance_4_L8), .Z(
        LED_128_Instance_subcells_out[18]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L4), .B(
        LED_128_Instance_SBox_Instance_4_T3), .Z(
        LED_128_Instance_subcells_out[17]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_4_L3), .B(
        LED_128_Instance_SBox_Instance_4_T2), .Z(
        LED_128_Instance_subcells_out[16]) );
  INV_X1 LED_128_Instance_SBox_Instance_5_U3 ( .A(
        LED_128_Instance_SBox_Instance_5_L0), .ZN(
        LED_128_Instance_SBox_Instance_5_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_5_U2 ( .A(
        LED_128_Instance_addconst_out[23]), .ZN(
        LED_128_Instance_SBox_Instance_5_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_5_U1 ( .A(
        LED_128_Instance_addconst_out[21]), .ZN(
        LED_128_Instance_SBox_Instance_5_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[22]), .B(
        LED_128_Instance_addconst_out[21]), .Z(
        LED_128_Instance_SBox_Instance_5_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[21]), .B(
        LED_128_Instance_addconst_out[20]), .Z(
        LED_128_Instance_SBox_Instance_5_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L1), .B(
        LED_128_Instance_addconst_out[23]), .Z(
        LED_128_Instance_SBox_Instance_5_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_T0), .B(
        LED_128_Instance_SBox_Instance_5_L2), .ZN(
        LED_128_Instance_SBox_Instance_5_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[23]), .B(
        LED_128_Instance_addconst_out[20]), .Z(
        LED_128_Instance_SBox_Instance_5_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L3), .B(
        LED_128_Instance_SBox_Instance_5_L0), .Z(
        LED_128_Instance_SBox_Instance_5_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[23]), .B(
        LED_128_Instance_addconst_out[21]), .Z(
        LED_128_Instance_SBox_Instance_5_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_T0), .B(
        LED_128_Instance_SBox_Instance_5_T2), .Z(
        LED_128_Instance_SBox_Instance_5_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L4), .B(
        LED_128_Instance_SBox_Instance_5_L5), .ZN(
        LED_128_Instance_SBox_Instance_5_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L1), .B(
        LED_128_Instance_addconst_out[22]), .Z(
        LED_128_Instance_SBox_Instance_5_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_5_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_5_n1), .A2(
        LED_128_Instance_SBox_Instance_5_n2), .ZN(
        LED_128_Instance_SBox_Instance_5_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_5_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_5_Q2), .A2(
        LED_128_Instance_SBox_Instance_5_Q3), .ZN(
        LED_128_Instance_SBox_Instance_5_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_5_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_5_n3), .A2(
        LED_128_Instance_addconst_out[22]), .ZN(
        LED_128_Instance_SBox_Instance_5_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_5_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_5_Q6), .A2(
        LED_128_Instance_SBox_Instance_5_Q7), .ZN(
        LED_128_Instance_SBox_Instance_5_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L5), .B(
        LED_128_Instance_SBox_Instance_5_T3), .Z(
        LED_128_Instance_SBox_Instance_5_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[20]), .B(
        LED_128_Instance_SBox_Instance_5_L7), .Z(
        LED_128_Instance_subcells_out[23]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L5), .B(
        LED_128_Instance_SBox_Instance_5_T1), .Z(
        LED_128_Instance_SBox_Instance_5_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L1), .B(
        LED_128_Instance_SBox_Instance_5_L8), .Z(
        LED_128_Instance_subcells_out[22]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L4), .B(
        LED_128_Instance_SBox_Instance_5_T3), .Z(
        LED_128_Instance_subcells_out[21]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_5_L3), .B(
        LED_128_Instance_SBox_Instance_5_T2), .Z(
        LED_128_Instance_subcells_out[20]) );
  INV_X1 LED_128_Instance_SBox_Instance_6_U3 ( .A(
        LED_128_Instance_SBox_Instance_6_L0), .ZN(
        LED_128_Instance_SBox_Instance_6_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_6_U2 ( .A(
        LED_128_Instance_addconst_out[27]), .ZN(
        LED_128_Instance_SBox_Instance_6_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_6_U1 ( .A(
        LED_128_Instance_addconst_out[25]), .ZN(
        LED_128_Instance_SBox_Instance_6_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[26]), .B(
        LED_128_Instance_addconst_out[25]), .Z(
        LED_128_Instance_SBox_Instance_6_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[25]), .B(
        LED_128_Instance_addconst_out[24]), .Z(
        LED_128_Instance_SBox_Instance_6_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L1), .B(
        LED_128_Instance_addconst_out[27]), .Z(
        LED_128_Instance_SBox_Instance_6_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_T0), .B(
        LED_128_Instance_SBox_Instance_6_L2), .ZN(
        LED_128_Instance_SBox_Instance_6_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[27]), .B(
        LED_128_Instance_addconst_out[24]), .Z(
        LED_128_Instance_SBox_Instance_6_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L3), .B(
        LED_128_Instance_SBox_Instance_6_L0), .Z(
        LED_128_Instance_SBox_Instance_6_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[27]), .B(
        LED_128_Instance_addconst_out[25]), .Z(
        LED_128_Instance_SBox_Instance_6_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_T0), .B(
        LED_128_Instance_SBox_Instance_6_T2), .Z(
        LED_128_Instance_SBox_Instance_6_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L4), .B(
        LED_128_Instance_SBox_Instance_6_L5), .ZN(
        LED_128_Instance_SBox_Instance_6_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L1), .B(
        LED_128_Instance_addconst_out[26]), .Z(
        LED_128_Instance_SBox_Instance_6_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_6_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_6_n1), .A2(
        LED_128_Instance_SBox_Instance_6_n2), .ZN(
        LED_128_Instance_SBox_Instance_6_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_6_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_6_Q2), .A2(
        LED_128_Instance_SBox_Instance_6_Q3), .ZN(
        LED_128_Instance_SBox_Instance_6_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_6_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_6_n3), .A2(
        LED_128_Instance_addconst_out[26]), .ZN(
        LED_128_Instance_SBox_Instance_6_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_6_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_6_Q6), .A2(
        LED_128_Instance_SBox_Instance_6_Q7), .ZN(
        LED_128_Instance_SBox_Instance_6_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L5), .B(
        LED_128_Instance_SBox_Instance_6_T3), .Z(
        LED_128_Instance_SBox_Instance_6_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[24]), .B(
        LED_128_Instance_SBox_Instance_6_L7), .Z(
        LED_128_Instance_subcells_out[27]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L5), .B(
        LED_128_Instance_SBox_Instance_6_T1), .Z(
        LED_128_Instance_SBox_Instance_6_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L1), .B(
        LED_128_Instance_SBox_Instance_6_L8), .Z(
        LED_128_Instance_subcells_out[26]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L4), .B(
        LED_128_Instance_SBox_Instance_6_T3), .Z(
        LED_128_Instance_subcells_out[25]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_6_L3), .B(
        LED_128_Instance_SBox_Instance_6_T2), .Z(
        LED_128_Instance_subcells_out[24]) );
  INV_X1 LED_128_Instance_SBox_Instance_7_U3 ( .A(
        LED_128_Instance_SBox_Instance_7_L0), .ZN(
        LED_128_Instance_SBox_Instance_7_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_7_U2 ( .A(
        LED_128_Instance_addconst_out[31]), .ZN(
        LED_128_Instance_SBox_Instance_7_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_7_U1 ( .A(
        LED_128_Instance_addconst_out[29]), .ZN(
        LED_128_Instance_SBox_Instance_7_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[30]), .B(
        LED_128_Instance_addconst_out[29]), .Z(
        LED_128_Instance_SBox_Instance_7_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[29]), .B(
        LED_128_Instance_addconst_out[28]), .Z(
        LED_128_Instance_SBox_Instance_7_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L1), .B(
        LED_128_Instance_addconst_out[31]), .Z(
        LED_128_Instance_SBox_Instance_7_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_T0), .B(
        LED_128_Instance_SBox_Instance_7_L2), .ZN(
        LED_128_Instance_SBox_Instance_7_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[31]), .B(
        LED_128_Instance_addconst_out[28]), .Z(
        LED_128_Instance_SBox_Instance_7_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L3), .B(
        LED_128_Instance_SBox_Instance_7_L0), .Z(
        LED_128_Instance_SBox_Instance_7_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[31]), .B(
        LED_128_Instance_addconst_out[29]), .Z(
        LED_128_Instance_SBox_Instance_7_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_T0), .B(
        LED_128_Instance_SBox_Instance_7_T2), .Z(
        LED_128_Instance_SBox_Instance_7_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L4), .B(
        LED_128_Instance_SBox_Instance_7_L5), .ZN(
        LED_128_Instance_SBox_Instance_7_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L1), .B(
        LED_128_Instance_addconst_out[30]), .Z(
        LED_128_Instance_SBox_Instance_7_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_7_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_7_n1), .A2(
        LED_128_Instance_SBox_Instance_7_n2), .ZN(
        LED_128_Instance_SBox_Instance_7_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_7_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_7_Q2), .A2(
        LED_128_Instance_SBox_Instance_7_Q3), .ZN(
        LED_128_Instance_SBox_Instance_7_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_7_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_7_n3), .A2(
        LED_128_Instance_addconst_out[30]), .ZN(
        LED_128_Instance_SBox_Instance_7_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_7_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_7_Q6), .A2(
        LED_128_Instance_SBox_Instance_7_Q7), .ZN(
        LED_128_Instance_SBox_Instance_7_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L5), .B(
        LED_128_Instance_SBox_Instance_7_T3), .Z(
        LED_128_Instance_SBox_Instance_7_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[28]), .B(
        LED_128_Instance_SBox_Instance_7_L7), .Z(
        LED_128_Instance_subcells_out[31]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L5), .B(
        LED_128_Instance_SBox_Instance_7_T1), .Z(
        LED_128_Instance_SBox_Instance_7_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L1), .B(
        LED_128_Instance_SBox_Instance_7_L8), .Z(
        LED_128_Instance_subcells_out[30]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L4), .B(
        LED_128_Instance_SBox_Instance_7_T3), .Z(
        LED_128_Instance_subcells_out[29]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_7_L3), .B(
        LED_128_Instance_SBox_Instance_7_T2), .Z(
        LED_128_Instance_subcells_out[28]) );
  INV_X1 LED_128_Instance_SBox_Instance_8_U3 ( .A(
        LED_128_Instance_SBox_Instance_8_L0), .ZN(
        LED_128_Instance_SBox_Instance_8_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_8_U2 ( .A(
        LED_128_Instance_addconst_out[35]), .ZN(
        LED_128_Instance_SBox_Instance_8_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_8_U1 ( .A(
        LED_128_Instance_addconst_out[33]), .ZN(
        LED_128_Instance_SBox_Instance_8_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[34]), .B(
        LED_128_Instance_addconst_out[33]), .Z(
        LED_128_Instance_SBox_Instance_8_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[33]), .B(
        LED_128_Instance_addconst_out[32]), .Z(
        LED_128_Instance_SBox_Instance_8_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L1), .B(
        LED_128_Instance_addconst_out[35]), .Z(
        LED_128_Instance_SBox_Instance_8_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_T0), .B(
        LED_128_Instance_SBox_Instance_8_L2), .ZN(
        LED_128_Instance_SBox_Instance_8_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[35]), .B(
        LED_128_Instance_addconst_out[32]), .Z(
        LED_128_Instance_SBox_Instance_8_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L3), .B(
        LED_128_Instance_SBox_Instance_8_L0), .Z(
        LED_128_Instance_SBox_Instance_8_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[35]), .B(
        LED_128_Instance_addconst_out[33]), .Z(
        LED_128_Instance_SBox_Instance_8_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_T0), .B(
        LED_128_Instance_SBox_Instance_8_T2), .Z(
        LED_128_Instance_SBox_Instance_8_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L4), .B(
        LED_128_Instance_SBox_Instance_8_L5), .ZN(
        LED_128_Instance_SBox_Instance_8_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L1), .B(
        LED_128_Instance_addconst_out[34]), .Z(
        LED_128_Instance_SBox_Instance_8_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_8_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_8_n1), .A2(
        LED_128_Instance_SBox_Instance_8_n2), .ZN(
        LED_128_Instance_SBox_Instance_8_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_8_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_8_Q2), .A2(
        LED_128_Instance_SBox_Instance_8_Q3), .ZN(
        LED_128_Instance_SBox_Instance_8_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_8_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_8_n3), .A2(
        LED_128_Instance_addconst_out[34]), .ZN(
        LED_128_Instance_SBox_Instance_8_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_8_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_8_Q6), .A2(
        LED_128_Instance_SBox_Instance_8_Q7), .ZN(
        LED_128_Instance_SBox_Instance_8_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L5), .B(
        LED_128_Instance_SBox_Instance_8_T3), .Z(
        LED_128_Instance_SBox_Instance_8_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[32]), .B(
        LED_128_Instance_SBox_Instance_8_L7), .Z(
        LED_128_Instance_subcells_out[35]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L5), .B(
        LED_128_Instance_SBox_Instance_8_T1), .Z(
        LED_128_Instance_SBox_Instance_8_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L1), .B(
        LED_128_Instance_SBox_Instance_8_L8), .Z(
        LED_128_Instance_subcells_out[34]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L4), .B(
        LED_128_Instance_SBox_Instance_8_T3), .Z(
        LED_128_Instance_subcells_out[33]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_8_L3), .B(
        LED_128_Instance_SBox_Instance_8_T2), .Z(
        LED_128_Instance_subcells_out[32]) );
  INV_X1 LED_128_Instance_SBox_Instance_9_U3 ( .A(
        LED_128_Instance_SBox_Instance_9_L0), .ZN(
        LED_128_Instance_SBox_Instance_9_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_9_U2 ( .A(
        LED_128_Instance_addconst_out[39]), .ZN(
        LED_128_Instance_SBox_Instance_9_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_9_U1 ( .A(
        LED_128_Instance_addconst_out[37]), .ZN(
        LED_128_Instance_SBox_Instance_9_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[38]), .B(
        LED_128_Instance_addconst_out[37]), .Z(
        LED_128_Instance_SBox_Instance_9_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[37]), .B(
        LED_128_Instance_addconst_out[36]), .Z(
        LED_128_Instance_SBox_Instance_9_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L1), .B(
        LED_128_Instance_addconst_out[39]), .Z(
        LED_128_Instance_SBox_Instance_9_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_T0), .B(
        LED_128_Instance_SBox_Instance_9_L2), .ZN(
        LED_128_Instance_SBox_Instance_9_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[39]), .B(
        LED_128_Instance_addconst_out[36]), .Z(
        LED_128_Instance_SBox_Instance_9_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L3), .B(
        LED_128_Instance_SBox_Instance_9_L0), .Z(
        LED_128_Instance_SBox_Instance_9_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[39]), .B(
        LED_128_Instance_addconst_out[37]), .Z(
        LED_128_Instance_SBox_Instance_9_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_T0), .B(
        LED_128_Instance_SBox_Instance_9_T2), .Z(
        LED_128_Instance_SBox_Instance_9_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L4), .B(
        LED_128_Instance_SBox_Instance_9_L5), .ZN(
        LED_128_Instance_SBox_Instance_9_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L1), .B(
        LED_128_Instance_addconst_out[38]), .Z(
        LED_128_Instance_SBox_Instance_9_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_9_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_9_n1), .A2(
        LED_128_Instance_SBox_Instance_9_n2), .ZN(
        LED_128_Instance_SBox_Instance_9_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_9_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_9_Q2), .A2(
        LED_128_Instance_SBox_Instance_9_Q3), .ZN(
        LED_128_Instance_SBox_Instance_9_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_9_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_9_n3), .A2(
        LED_128_Instance_addconst_out[38]), .ZN(
        LED_128_Instance_SBox_Instance_9_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_9_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_9_Q6), .A2(
        LED_128_Instance_SBox_Instance_9_Q7), .ZN(
        LED_128_Instance_SBox_Instance_9_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L5), .B(
        LED_128_Instance_SBox_Instance_9_T3), .Z(
        LED_128_Instance_SBox_Instance_9_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[36]), .B(
        LED_128_Instance_SBox_Instance_9_L7), .Z(
        LED_128_Instance_subcells_out[39]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L5), .B(
        LED_128_Instance_SBox_Instance_9_T1), .Z(
        LED_128_Instance_SBox_Instance_9_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L1), .B(
        LED_128_Instance_SBox_Instance_9_L8), .Z(
        LED_128_Instance_subcells_out[38]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L4), .B(
        LED_128_Instance_SBox_Instance_9_T3), .Z(
        LED_128_Instance_subcells_out[37]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_9_L3), .B(
        LED_128_Instance_SBox_Instance_9_T2), .Z(
        LED_128_Instance_subcells_out[36]) );
  INV_X1 LED_128_Instance_SBox_Instance_10_U3 ( .A(
        LED_128_Instance_SBox_Instance_10_L0), .ZN(
        LED_128_Instance_SBox_Instance_10_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_10_U2 ( .A(
        LED_128_Instance_addconst_out[43]), .ZN(
        LED_128_Instance_SBox_Instance_10_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_10_U1 ( .A(
        LED_128_Instance_addconst_out[41]), .ZN(
        LED_128_Instance_SBox_Instance_10_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[42]), .B(
        LED_128_Instance_addconst_out[41]), .Z(
        LED_128_Instance_SBox_Instance_10_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[41]), .B(
        LED_128_Instance_addconst_out[40]), .Z(
        LED_128_Instance_SBox_Instance_10_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L1), .B(
        LED_128_Instance_addconst_out[43]), .Z(
        LED_128_Instance_SBox_Instance_10_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_T0), .B(
        LED_128_Instance_SBox_Instance_10_L2), .ZN(
        LED_128_Instance_SBox_Instance_10_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[43]), .B(
        LED_128_Instance_addconst_out[40]), .Z(
        LED_128_Instance_SBox_Instance_10_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L3), .B(
        LED_128_Instance_SBox_Instance_10_L0), .Z(
        LED_128_Instance_SBox_Instance_10_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[43]), .B(
        LED_128_Instance_addconst_out[41]), .Z(
        LED_128_Instance_SBox_Instance_10_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_T0), .B(
        LED_128_Instance_SBox_Instance_10_T2), .Z(
        LED_128_Instance_SBox_Instance_10_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L4), .B(
        LED_128_Instance_SBox_Instance_10_L5), .ZN(
        LED_128_Instance_SBox_Instance_10_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L1), .B(
        LED_128_Instance_addconst_out[42]), .Z(
        LED_128_Instance_SBox_Instance_10_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_10_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_10_n1), .A2(
        LED_128_Instance_SBox_Instance_10_n2), .ZN(
        LED_128_Instance_SBox_Instance_10_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_10_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_10_Q2), .A2(
        LED_128_Instance_SBox_Instance_10_Q3), .ZN(
        LED_128_Instance_SBox_Instance_10_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_10_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_10_n3), .A2(
        LED_128_Instance_addconst_out[42]), .ZN(
        LED_128_Instance_SBox_Instance_10_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_10_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_10_Q6), .A2(
        LED_128_Instance_SBox_Instance_10_Q7), .ZN(
        LED_128_Instance_SBox_Instance_10_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L5), .B(
        LED_128_Instance_SBox_Instance_10_T3), .Z(
        LED_128_Instance_SBox_Instance_10_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[40]), .B(
        LED_128_Instance_SBox_Instance_10_L7), .Z(
        LED_128_Instance_subcells_out[43]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L5), .B(
        LED_128_Instance_SBox_Instance_10_T1), .Z(
        LED_128_Instance_SBox_Instance_10_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L1), .B(
        LED_128_Instance_SBox_Instance_10_L8), .Z(
        LED_128_Instance_subcells_out[42]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L4), .B(
        LED_128_Instance_SBox_Instance_10_T3), .Z(
        LED_128_Instance_subcells_out[41]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_10_L3), .B(
        LED_128_Instance_SBox_Instance_10_T2), .Z(
        LED_128_Instance_subcells_out[40]) );
  INV_X1 LED_128_Instance_SBox_Instance_11_U3 ( .A(
        LED_128_Instance_SBox_Instance_11_L0), .ZN(
        LED_128_Instance_SBox_Instance_11_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_11_U2 ( .A(
        LED_128_Instance_addconst_out[47]), .ZN(
        LED_128_Instance_SBox_Instance_11_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_11_U1 ( .A(
        LED_128_Instance_addconst_out[45]), .ZN(
        LED_128_Instance_SBox_Instance_11_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[46]), .B(
        LED_128_Instance_addconst_out[45]), .Z(
        LED_128_Instance_SBox_Instance_11_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[45]), .B(
        LED_128_Instance_addconst_out[44]), .Z(
        LED_128_Instance_SBox_Instance_11_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L1), .B(
        LED_128_Instance_addconst_out[47]), .Z(
        LED_128_Instance_SBox_Instance_11_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_T0), .B(
        LED_128_Instance_SBox_Instance_11_L2), .ZN(
        LED_128_Instance_SBox_Instance_11_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[47]), .B(
        LED_128_Instance_addconst_out[44]), .Z(
        LED_128_Instance_SBox_Instance_11_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L3), .B(
        LED_128_Instance_SBox_Instance_11_L0), .Z(
        LED_128_Instance_SBox_Instance_11_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[47]), .B(
        LED_128_Instance_addconst_out[45]), .Z(
        LED_128_Instance_SBox_Instance_11_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_T0), .B(
        LED_128_Instance_SBox_Instance_11_T2), .Z(
        LED_128_Instance_SBox_Instance_11_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L4), .B(
        LED_128_Instance_SBox_Instance_11_L5), .ZN(
        LED_128_Instance_SBox_Instance_11_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L1), .B(
        LED_128_Instance_addconst_out[46]), .Z(
        LED_128_Instance_SBox_Instance_11_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_11_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_11_n1), .A2(
        LED_128_Instance_SBox_Instance_11_n2), .ZN(
        LED_128_Instance_SBox_Instance_11_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_11_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_11_Q2), .A2(
        LED_128_Instance_SBox_Instance_11_Q3), .ZN(
        LED_128_Instance_SBox_Instance_11_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_11_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_11_n3), .A2(
        LED_128_Instance_addconst_out[46]), .ZN(
        LED_128_Instance_SBox_Instance_11_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_11_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_11_Q6), .A2(
        LED_128_Instance_SBox_Instance_11_Q7), .ZN(
        LED_128_Instance_SBox_Instance_11_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L5), .B(
        LED_128_Instance_SBox_Instance_11_T3), .Z(
        LED_128_Instance_SBox_Instance_11_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[44]), .B(
        LED_128_Instance_SBox_Instance_11_L7), .Z(
        LED_128_Instance_subcells_out[47]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L5), .B(
        LED_128_Instance_SBox_Instance_11_T1), .Z(
        LED_128_Instance_SBox_Instance_11_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L1), .B(
        LED_128_Instance_SBox_Instance_11_L8), .Z(
        LED_128_Instance_subcells_out[46]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L4), .B(
        LED_128_Instance_SBox_Instance_11_T3), .Z(
        LED_128_Instance_subcells_out[45]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_11_L3), .B(
        LED_128_Instance_SBox_Instance_11_T2), .Z(
        LED_128_Instance_subcells_out[44]) );
  INV_X1 LED_128_Instance_SBox_Instance_12_U3 ( .A(
        LED_128_Instance_SBox_Instance_12_L0), .ZN(
        LED_128_Instance_SBox_Instance_12_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_12_U2 ( .A(
        LED_128_Instance_addconst_out[51]), .ZN(
        LED_128_Instance_SBox_Instance_12_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_12_U1 ( .A(
        LED_128_Instance_addconst_out[49]), .ZN(
        LED_128_Instance_SBox_Instance_12_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[50]), .B(
        LED_128_Instance_addconst_out[49]), .Z(
        LED_128_Instance_SBox_Instance_12_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[49]), .B(
        LED_128_Instance_addconst_out[48]), .Z(
        LED_128_Instance_SBox_Instance_12_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L1), .B(
        LED_128_Instance_addconst_out[51]), .Z(
        LED_128_Instance_SBox_Instance_12_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_T0), .B(
        LED_128_Instance_SBox_Instance_12_L2), .ZN(
        LED_128_Instance_SBox_Instance_12_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[51]), .B(
        LED_128_Instance_addconst_out[48]), .Z(
        LED_128_Instance_SBox_Instance_12_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L3), .B(
        LED_128_Instance_SBox_Instance_12_L0), .Z(
        LED_128_Instance_SBox_Instance_12_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[51]), .B(
        LED_128_Instance_addconst_out[49]), .Z(
        LED_128_Instance_SBox_Instance_12_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_T0), .B(
        LED_128_Instance_SBox_Instance_12_T2), .Z(
        LED_128_Instance_SBox_Instance_12_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L4), .B(
        LED_128_Instance_SBox_Instance_12_L5), .ZN(
        LED_128_Instance_SBox_Instance_12_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L1), .B(
        LED_128_Instance_addconst_out[50]), .Z(
        LED_128_Instance_SBox_Instance_12_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_12_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_12_n1), .A2(
        LED_128_Instance_SBox_Instance_12_n2), .ZN(
        LED_128_Instance_SBox_Instance_12_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_12_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_12_Q2), .A2(
        LED_128_Instance_SBox_Instance_12_Q3), .ZN(
        LED_128_Instance_SBox_Instance_12_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_12_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_12_n3), .A2(
        LED_128_Instance_addconst_out[50]), .ZN(
        LED_128_Instance_SBox_Instance_12_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_12_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_12_Q6), .A2(
        LED_128_Instance_SBox_Instance_12_Q7), .ZN(
        LED_128_Instance_SBox_Instance_12_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L5), .B(
        LED_128_Instance_SBox_Instance_12_T3), .Z(
        LED_128_Instance_SBox_Instance_12_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[48]), .B(
        LED_128_Instance_SBox_Instance_12_L7), .Z(
        LED_128_Instance_subcells_out[51]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L5), .B(
        LED_128_Instance_SBox_Instance_12_T1), .Z(
        LED_128_Instance_SBox_Instance_12_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L1), .B(
        LED_128_Instance_SBox_Instance_12_L8), .Z(
        LED_128_Instance_subcells_out[50]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L4), .B(
        LED_128_Instance_SBox_Instance_12_T3), .Z(
        LED_128_Instance_subcells_out[49]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_12_L3), .B(
        LED_128_Instance_SBox_Instance_12_T2), .Z(
        LED_128_Instance_subcells_out[48]) );
  INV_X1 LED_128_Instance_SBox_Instance_13_U3 ( .A(
        LED_128_Instance_SBox_Instance_13_L0), .ZN(
        LED_128_Instance_SBox_Instance_13_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_13_U2 ( .A(
        LED_128_Instance_addconst_out[55]), .ZN(
        LED_128_Instance_SBox_Instance_13_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_13_U1 ( .A(
        LED_128_Instance_addconst_out[53]), .ZN(
        LED_128_Instance_SBox_Instance_13_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[54]), .B(
        LED_128_Instance_addconst_out[53]), .Z(
        LED_128_Instance_SBox_Instance_13_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[53]), .B(
        LED_128_Instance_addconst_out[52]), .Z(
        LED_128_Instance_SBox_Instance_13_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L1), .B(
        LED_128_Instance_addconst_out[55]), .Z(
        LED_128_Instance_SBox_Instance_13_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_T0), .B(
        LED_128_Instance_SBox_Instance_13_L2), .ZN(
        LED_128_Instance_SBox_Instance_13_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[55]), .B(
        LED_128_Instance_addconst_out[52]), .Z(
        LED_128_Instance_SBox_Instance_13_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L3), .B(
        LED_128_Instance_SBox_Instance_13_L0), .Z(
        LED_128_Instance_SBox_Instance_13_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[55]), .B(
        LED_128_Instance_addconst_out[53]), .Z(
        LED_128_Instance_SBox_Instance_13_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_T0), .B(
        LED_128_Instance_SBox_Instance_13_T2), .Z(
        LED_128_Instance_SBox_Instance_13_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L4), .B(
        LED_128_Instance_SBox_Instance_13_L5), .ZN(
        LED_128_Instance_SBox_Instance_13_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L1), .B(
        LED_128_Instance_addconst_out[54]), .Z(
        LED_128_Instance_SBox_Instance_13_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_13_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_13_n1), .A2(
        LED_128_Instance_SBox_Instance_13_n2), .ZN(
        LED_128_Instance_SBox_Instance_13_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_13_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_13_Q2), .A2(
        LED_128_Instance_SBox_Instance_13_Q3), .ZN(
        LED_128_Instance_SBox_Instance_13_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_13_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_13_n3), .A2(
        LED_128_Instance_addconst_out[54]), .ZN(
        LED_128_Instance_SBox_Instance_13_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_13_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_13_Q6), .A2(
        LED_128_Instance_SBox_Instance_13_Q7), .ZN(
        LED_128_Instance_SBox_Instance_13_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L5), .B(
        LED_128_Instance_SBox_Instance_13_T3), .Z(
        LED_128_Instance_SBox_Instance_13_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[52]), .B(
        LED_128_Instance_SBox_Instance_13_L7), .Z(
        LED_128_Instance_subcells_out[55]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L5), .B(
        LED_128_Instance_SBox_Instance_13_T1), .Z(
        LED_128_Instance_SBox_Instance_13_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L1), .B(
        LED_128_Instance_SBox_Instance_13_L8), .Z(
        LED_128_Instance_subcells_out[54]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L4), .B(
        LED_128_Instance_SBox_Instance_13_T3), .Z(
        LED_128_Instance_subcells_out[53]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_13_L3), .B(
        LED_128_Instance_SBox_Instance_13_T2), .Z(
        LED_128_Instance_subcells_out[52]) );
  INV_X1 LED_128_Instance_SBox_Instance_14_U3 ( .A(
        LED_128_Instance_SBox_Instance_14_L0), .ZN(
        LED_128_Instance_SBox_Instance_14_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_14_U2 ( .A(
        LED_128_Instance_addconst_out[59]), .ZN(
        LED_128_Instance_SBox_Instance_14_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_14_U1 ( .A(
        LED_128_Instance_addconst_out[57]), .ZN(
        LED_128_Instance_SBox_Instance_14_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[58]), .B(
        LED_128_Instance_addconst_out[57]), .Z(
        LED_128_Instance_SBox_Instance_14_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[57]), .B(
        LED_128_Instance_addconst_out[56]), .Z(
        LED_128_Instance_SBox_Instance_14_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L1), .B(
        LED_128_Instance_addconst_out[59]), .Z(
        LED_128_Instance_SBox_Instance_14_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_T0), .B(
        LED_128_Instance_SBox_Instance_14_L2), .ZN(
        LED_128_Instance_SBox_Instance_14_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[59]), .B(
        LED_128_Instance_addconst_out[56]), .Z(
        LED_128_Instance_SBox_Instance_14_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L3), .B(
        LED_128_Instance_SBox_Instance_14_L0), .Z(
        LED_128_Instance_SBox_Instance_14_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[59]), .B(
        LED_128_Instance_addconst_out[57]), .Z(
        LED_128_Instance_SBox_Instance_14_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_T0), .B(
        LED_128_Instance_SBox_Instance_14_T2), .Z(
        LED_128_Instance_SBox_Instance_14_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L4), .B(
        LED_128_Instance_SBox_Instance_14_L5), .ZN(
        LED_128_Instance_SBox_Instance_14_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L1), .B(
        LED_128_Instance_addconst_out[58]), .Z(
        LED_128_Instance_SBox_Instance_14_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_14_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_14_n1), .A2(
        LED_128_Instance_SBox_Instance_14_n2), .ZN(
        LED_128_Instance_SBox_Instance_14_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_14_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_14_Q2), .A2(
        LED_128_Instance_SBox_Instance_14_Q3), .ZN(
        LED_128_Instance_SBox_Instance_14_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_14_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_14_n3), .A2(
        LED_128_Instance_addconst_out[58]), .ZN(
        LED_128_Instance_SBox_Instance_14_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_14_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_14_Q6), .A2(
        LED_128_Instance_SBox_Instance_14_Q7), .ZN(
        LED_128_Instance_SBox_Instance_14_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L5), .B(
        LED_128_Instance_SBox_Instance_14_T3), .Z(
        LED_128_Instance_SBox_Instance_14_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[56]), .B(
        LED_128_Instance_SBox_Instance_14_L7), .Z(
        LED_128_Instance_subcells_out[59]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L5), .B(
        LED_128_Instance_SBox_Instance_14_T1), .Z(
        LED_128_Instance_SBox_Instance_14_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L1), .B(
        LED_128_Instance_SBox_Instance_14_L8), .Z(
        LED_128_Instance_subcells_out[58]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L4), .B(
        LED_128_Instance_SBox_Instance_14_T3), .Z(
        LED_128_Instance_subcells_out[57]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_14_L3), .B(
        LED_128_Instance_SBox_Instance_14_T2), .Z(
        LED_128_Instance_subcells_out[56]) );
  INV_X1 LED_128_Instance_SBox_Instance_15_U3 ( .A(
        LED_128_Instance_SBox_Instance_15_L0), .ZN(
        LED_128_Instance_SBox_Instance_15_n1) );
  INV_X1 LED_128_Instance_SBox_Instance_15_U2 ( .A(
        LED_128_Instance_addconst_out[63]), .ZN(
        LED_128_Instance_SBox_Instance_15_n2) );
  INV_X1 LED_128_Instance_SBox_Instance_15_U1 ( .A(
        LED_128_Instance_addconst_out[61]), .ZN(
        LED_128_Instance_SBox_Instance_15_n3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .A(
        LED_128_Instance_addconst_out[62]), .B(
        LED_128_Instance_addconst_out[61]), .Z(
        LED_128_Instance_SBox_Instance_15_L0) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .A(
        LED_128_Instance_addconst_out[61]), .B(
        LED_128_Instance_addconst_out[60]), .Z(
        LED_128_Instance_SBox_Instance_15_L1) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L1), .B(
        LED_128_Instance_addconst_out[63]), .Z(
        LED_128_Instance_SBox_Instance_15_L2) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_T0), .B(
        LED_128_Instance_SBox_Instance_15_L2), .ZN(
        LED_128_Instance_SBox_Instance_15_Q2) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .A(
        LED_128_Instance_addconst_out[63]), .B(
        LED_128_Instance_addconst_out[60]), .Z(
        LED_128_Instance_SBox_Instance_15_L3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L3), .B(
        LED_128_Instance_SBox_Instance_15_L0), .Z(
        LED_128_Instance_SBox_Instance_15_Q3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .A(
        LED_128_Instance_addconst_out[63]), .B(
        LED_128_Instance_addconst_out[61]), .Z(
        LED_128_Instance_SBox_Instance_15_L4) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_T0), .B(
        LED_128_Instance_SBox_Instance_15_T2), .Z(
        LED_128_Instance_SBox_Instance_15_L5) );
  XNOR2_X1 LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L4), .B(
        LED_128_Instance_SBox_Instance_15_L5), .ZN(
        LED_128_Instance_SBox_Instance_15_Q6) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L1), .B(
        LED_128_Instance_addconst_out[62]), .Z(
        LED_128_Instance_SBox_Instance_15_Q7) );
  AND2_X1 LED_128_Instance_SBox_Instance_15_AND1_U1 ( .A1(
        LED_128_Instance_SBox_Instance_15_n1), .A2(
        LED_128_Instance_SBox_Instance_15_n2), .ZN(
        LED_128_Instance_SBox_Instance_15_T0) );
  AND2_X1 LED_128_Instance_SBox_Instance_15_AND2_U1 ( .A1(
        LED_128_Instance_SBox_Instance_15_Q2), .A2(
        LED_128_Instance_SBox_Instance_15_Q3), .ZN(
        LED_128_Instance_SBox_Instance_15_T1) );
  AND2_X1 LED_128_Instance_SBox_Instance_15_AND3_U1 ( .A1(
        LED_128_Instance_SBox_Instance_15_n3), .A2(
        LED_128_Instance_addconst_out[62]), .ZN(
        LED_128_Instance_SBox_Instance_15_T2) );
  AND2_X1 LED_128_Instance_SBox_Instance_15_AND4_U1 ( .A1(
        LED_128_Instance_SBox_Instance_15_Q6), .A2(
        LED_128_Instance_SBox_Instance_15_Q7), .ZN(
        LED_128_Instance_SBox_Instance_15_T3) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L5), .B(
        LED_128_Instance_SBox_Instance_15_T3), .Z(
        LED_128_Instance_SBox_Instance_15_L7) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .A(
        LED_128_Instance_addconst_out[60]), .B(
        LED_128_Instance_SBox_Instance_15_L7), .Z(
        LED_128_Instance_subcells_out[63]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L5), .B(
        LED_128_Instance_SBox_Instance_15_T1), .Z(
        LED_128_Instance_SBox_Instance_15_L8) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L1), .B(
        LED_128_Instance_SBox_Instance_15_L8), .Z(
        LED_128_Instance_subcells_out[62]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L4), .B(
        LED_128_Instance_SBox_Instance_15_T3), .Z(
        LED_128_Instance_subcells_out[61]) );
  XOR2_X1 LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .A(
        LED_128_Instance_SBox_Instance_15_L3), .B(
        LED_128_Instance_SBox_Instance_15_T2), .Z(
        LED_128_Instance_subcells_out[60]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U54 ( .A(
        LED_128_Instance_MCS_Instance_0_n38), .B(
        LED_128_Instance_MCS_Instance_0_n37), .ZN(
        LED_128_Instance_mixcolumns_out[51]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U53 ( .A(
        LED_128_Instance_mixcolumns_out[3]), .B(
        LED_128_Instance_subcells_out[61]), .ZN(
        LED_128_Instance_MCS_Instance_0_n37) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U52 ( .A(
        LED_128_Instance_mixcolumns_out[34]), .B(
        LED_128_Instance_mixcolumns_out[18]), .Z(
        LED_128_Instance_MCS_Instance_0_n38) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U51 ( .A(
        LED_128_Instance_MCS_Instance_0_n36), .B(
        LED_128_Instance_MCS_Instance_0_n35), .ZN(
        LED_128_Instance_mixcolumns_out[34]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U50 ( .A(
        LED_128_Instance_subcells_out[62]), .B(
        LED_128_Instance_MCS_Instance_0_n34), .ZN(
        LED_128_Instance_MCS_Instance_0_n36) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U49 ( .A(
        LED_128_Instance_MCS_Instance_0_n33), .B(
        LED_128_Instance_mixcolumns_out[33]), .ZN(
        LED_128_Instance_mixcolumns_out[50]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U48 ( .A(
        LED_128_Instance_mixcolumns_out[2]), .B(
        LED_128_Instance_MCS_Instance_0_n35), .ZN(
        LED_128_Instance_MCS_Instance_0_n33) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U47 ( .A(
        LED_128_Instance_MCS_Instance_0_n32), .B(
        LED_128_Instance_MCS_Instance_0_n31), .ZN(
        LED_128_Instance_mixcolumns_out[49]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U46 ( .A(
        LED_128_Instance_MCS_Instance_0_n30), .B(
        LED_128_Instance_MCS_Instance_0_n29), .ZN(
        LED_128_Instance_MCS_Instance_0_n32) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U45 ( .A(
        LED_128_Instance_subcells_out[63]), .B(
        LED_128_Instance_mixcolumns_out[1]), .ZN(
        LED_128_Instance_MCS_Instance_0_n29) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U44 ( .A(
        LED_128_Instance_mixcolumns_out[32]), .B(
        LED_128_Instance_MCS_Instance_0_n28), .Z(
        LED_128_Instance_MCS_Instance_0_n30) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U43 ( .A(
        LED_128_Instance_MCS_Instance_0_n27), .B(
        LED_128_Instance_MCS_Instance_0_n26), .ZN(
        LED_128_Instance_mixcolumns_out[32]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U42 ( .A(
        LED_128_Instance_subcells_out[42]), .B(
        LED_128_Instance_mixcolumns_out[3]), .ZN(
        LED_128_Instance_MCS_Instance_0_n26) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U41 ( .A(
        LED_128_Instance_subcells_out[60]), .B(
        LED_128_Instance_mixcolumns_out[19]), .Z(
        LED_128_Instance_MCS_Instance_0_n27) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U40 ( .A(
        LED_128_Instance_MCS_Instance_0_n25), .B(
        LED_128_Instance_mixcolumns_out[0]), .ZN(
        LED_128_Instance_mixcolumns_out[48]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U39 ( .A(
        LED_128_Instance_mixcolumns_out[19]), .B(
        LED_128_Instance_MCS_Instance_0_n28), .ZN(
        LED_128_Instance_MCS_Instance_0_n25) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U38 ( .A(
        LED_128_Instance_subcells_out[62]), .B(
        LED_128_Instance_mixcolumns_out[35]), .Z(
        LED_128_Instance_MCS_Instance_0_n28) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U37 ( .A(
        LED_128_Instance_MCS_Instance_0_n24), .B(
        LED_128_Instance_MCS_Instance_0_n23), .ZN(
        LED_128_Instance_mixcolumns_out[35]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U36 ( .A(
        LED_128_Instance_subcells_out[63]), .B(
        LED_128_Instance_subcells_out[41]), .ZN(
        LED_128_Instance_MCS_Instance_0_n23) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U35 ( .A(
        LED_128_Instance_mixcolumns_out[18]), .B(
        LED_128_Instance_mixcolumns_out[2]), .Z(
        LED_128_Instance_MCS_Instance_0_n24) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U34 ( .A(
        LED_128_Instance_MCS_Instance_0_n22), .B(
        LED_128_Instance_MCS_Instance_0_n21), .ZN(
        LED_128_Instance_mixcolumns_out[18]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U33 ( .A(
        LED_128_Instance_MCS_Instance_0_n20), .B(
        LED_128_Instance_subcells_out[61]), .ZN(
        LED_128_Instance_MCS_Instance_0_n21) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U32 ( .A(
        LED_128_Instance_mixcolumns_out[1]), .B(
        LED_128_Instance_subcells_out[20]), .Z(
        LED_128_Instance_MCS_Instance_0_n22) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U31 ( .A(
        LED_128_Instance_MCS_Instance_0_n19), .B(
        LED_128_Instance_MCS_Instance_0_n18), .ZN(
        LED_128_Instance_mixcolumns_out[1]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U30 ( .A(
        LED_128_Instance_subcells_out[40]), .B(
        LED_128_Instance_subcells_out[43]), .ZN(
        LED_128_Instance_MCS_Instance_0_n18) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U29 ( .A(
        LED_128_Instance_MCS_Instance_0_n17), .B(
        LED_128_Instance_MCS_Instance_0_n34), .Z(
        LED_128_Instance_MCS_Instance_0_n19) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U28 ( .A(
        LED_128_Instance_MCS_Instance_0_n16), .B(
        LED_128_Instance_subcells_out[2]), .ZN(
        LED_128_Instance_MCS_Instance_0_n34) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U27 ( .A(
        LED_128_Instance_subcells_out[21]), .B(
        LED_128_Instance_subcells_out[3]), .ZN(
        LED_128_Instance_MCS_Instance_0_n16) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U26 ( .A(
        LED_128_Instance_MCS_Instance_0_n15), .B(
        LED_128_Instance_MCS_Instance_0_n31), .ZN(
        LED_128_Instance_mixcolumns_out[33]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U25 ( .A(
        LED_128_Instance_mixcolumns_out[16]), .B(
        LED_128_Instance_mixcolumns_out[19]), .ZN(
        LED_128_Instance_MCS_Instance_0_n31) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U24 ( .A(
        LED_128_Instance_MCS_Instance_0_n14), .B(
        LED_128_Instance_MCS_Instance_0_n13), .ZN(
        LED_128_Instance_MCS_Instance_0_n15) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U23 ( .A(
        LED_128_Instance_subcells_out[42]), .B(
        LED_128_Instance_subcells_out[43]), .ZN(
        LED_128_Instance_MCS_Instance_0_n13) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U22 ( .A(
        LED_128_Instance_MCS_Instance_0_n12), .B(
        LED_128_Instance_subcells_out[61]), .Z(
        LED_128_Instance_MCS_Instance_0_n14) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U21 ( .A(
        LED_128_Instance_MCS_Instance_0_n11), .B(
        LED_128_Instance_MCS_Instance_0_n10), .ZN(
        LED_128_Instance_mixcolumns_out[16]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U20 ( .A(
        LED_128_Instance_mixcolumns_out[3]), .B(
        LED_128_Instance_subcells_out[63]), .ZN(
        LED_128_Instance_MCS_Instance_0_n10) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U19 ( .A(
        LED_128_Instance_subcells_out[40]), .B(
        LED_128_Instance_subcells_out[22]), .Z(
        LED_128_Instance_MCS_Instance_0_n11) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U18 ( .A(
        LED_128_Instance_MCS_Instance_0_n9), .B(
        LED_128_Instance_MCS_Instance_0_n8), .ZN(
        LED_128_Instance_mixcolumns_out[19]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U17 ( .A(
        LED_128_Instance_subcells_out[62]), .B(
        LED_128_Instance_subcells_out[43]), .ZN(
        LED_128_Instance_MCS_Instance_0_n8) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U16 ( .A(
        LED_128_Instance_mixcolumns_out[2]), .B(
        LED_128_Instance_subcells_out[21]), .Z(
        LED_128_Instance_MCS_Instance_0_n9) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U15 ( .A(
        LED_128_Instance_MCS_Instance_0_n7), .B(
        LED_128_Instance_MCS_Instance_0_n6), .ZN(
        LED_128_Instance_mixcolumns_out[2]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U14 ( .A(
        LED_128_Instance_MCS_Instance_0_n5), .B(
        LED_128_Instance_subcells_out[3]), .ZN(
        LED_128_Instance_MCS_Instance_0_n6) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U13 ( .A(
        LED_128_Instance_subcells_out[0]), .B(
        LED_128_Instance_subcells_out[61]), .Z(
        LED_128_Instance_MCS_Instance_0_n7) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U12 ( .A(
        LED_128_Instance_MCS_Instance_0_n17), .B(
        LED_128_Instance_MCS_Instance_0_n35), .Z(
        LED_128_Instance_mixcolumns_out[17]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U11 ( .A(
        LED_128_Instance_MCS_Instance_0_n4), .B(
        LED_128_Instance_MCS_Instance_0_n12), .ZN(
        LED_128_Instance_MCS_Instance_0_n35) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U10 ( .A(
        LED_128_Instance_mixcolumns_out[3]), .B(
        LED_128_Instance_mixcolumns_out[0]), .Z(
        LED_128_Instance_MCS_Instance_0_n12) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U9 ( .A(
        LED_128_Instance_subcells_out[23]), .B(
        LED_128_Instance_MCS_Instance_0_n5), .ZN(
        LED_128_Instance_MCS_Instance_0_n4) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U8 ( .A(
        LED_128_Instance_subcells_out[22]), .B(
        LED_128_Instance_subcells_out[41]), .Z(
        LED_128_Instance_MCS_Instance_0_n5) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U7 ( .A(
        LED_128_Instance_subcells_out[63]), .B(
        LED_128_Instance_subcells_out[60]), .Z(
        LED_128_Instance_MCS_Instance_0_n17) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U6 ( .A(
        LED_128_Instance_MCS_Instance_0_n3), .B(
        LED_128_Instance_MCS_Instance_0_n2), .ZN(
        LED_128_Instance_mixcolumns_out[0]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U5 ( .A(
        LED_128_Instance_subcells_out[63]), .B(
        LED_128_Instance_subcells_out[43]), .ZN(
        LED_128_Instance_MCS_Instance_0_n2) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U4 ( .A(
        LED_128_Instance_subcells_out[2]), .B(
        LED_128_Instance_subcells_out[20]), .Z(
        LED_128_Instance_MCS_Instance_0_n3) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U3 ( .A(
        LED_128_Instance_MCS_Instance_0_n1), .B(
        LED_128_Instance_subcells_out[62]), .ZN(
        LED_128_Instance_mixcolumns_out[3]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_0_U2 ( .A(
        LED_128_Instance_MCS_Instance_0_n20), .B(
        LED_128_Instance_subcells_out[1]), .ZN(
        LED_128_Instance_MCS_Instance_0_n1) );
  XOR2_X1 LED_128_Instance_MCS_Instance_0_U1 ( .A(
        LED_128_Instance_subcells_out[42]), .B(
        LED_128_Instance_subcells_out[23]), .Z(
        LED_128_Instance_MCS_Instance_0_n20) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U54 ( .A(
        LED_128_Instance_MCS_Instance_1_n38), .B(
        LED_128_Instance_MCS_Instance_1_n37), .ZN(
        LED_128_Instance_mixcolumns_out[55]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U53 ( .A(
        LED_128_Instance_mixcolumns_out[7]), .B(
        LED_128_Instance_subcells_out[49]), .ZN(
        LED_128_Instance_MCS_Instance_1_n37) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U52 ( .A(
        LED_128_Instance_mixcolumns_out[38]), .B(
        LED_128_Instance_mixcolumns_out[22]), .Z(
        LED_128_Instance_MCS_Instance_1_n38) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U51 ( .A(
        LED_128_Instance_MCS_Instance_1_n36), .B(
        LED_128_Instance_MCS_Instance_1_n35), .ZN(
        LED_128_Instance_mixcolumns_out[38]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U50 ( .A(
        LED_128_Instance_subcells_out[50]), .B(
        LED_128_Instance_MCS_Instance_1_n34), .ZN(
        LED_128_Instance_MCS_Instance_1_n36) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U49 ( .A(
        LED_128_Instance_MCS_Instance_1_n33), .B(
        LED_128_Instance_mixcolumns_out[37]), .ZN(
        LED_128_Instance_mixcolumns_out[54]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U48 ( .A(
        LED_128_Instance_mixcolumns_out[6]), .B(
        LED_128_Instance_MCS_Instance_1_n35), .ZN(
        LED_128_Instance_MCS_Instance_1_n33) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U47 ( .A(
        LED_128_Instance_MCS_Instance_1_n32), .B(
        LED_128_Instance_MCS_Instance_1_n31), .ZN(
        LED_128_Instance_mixcolumns_out[53]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U46 ( .A(
        LED_128_Instance_MCS_Instance_1_n30), .B(
        LED_128_Instance_MCS_Instance_1_n29), .ZN(
        LED_128_Instance_MCS_Instance_1_n32) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U45 ( .A(
        LED_128_Instance_subcells_out[51]), .B(
        LED_128_Instance_mixcolumns_out[5]), .ZN(
        LED_128_Instance_MCS_Instance_1_n29) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U44 ( .A(
        LED_128_Instance_mixcolumns_out[36]), .B(
        LED_128_Instance_MCS_Instance_1_n28), .Z(
        LED_128_Instance_MCS_Instance_1_n30) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U43 ( .A(
        LED_128_Instance_MCS_Instance_1_n27), .B(
        LED_128_Instance_MCS_Instance_1_n26), .ZN(
        LED_128_Instance_mixcolumns_out[36]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U42 ( .A(
        LED_128_Instance_subcells_out[46]), .B(
        LED_128_Instance_mixcolumns_out[7]), .ZN(
        LED_128_Instance_MCS_Instance_1_n26) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U41 ( .A(
        LED_128_Instance_subcells_out[48]), .B(
        LED_128_Instance_mixcolumns_out[23]), .Z(
        LED_128_Instance_MCS_Instance_1_n27) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U40 ( .A(
        LED_128_Instance_MCS_Instance_1_n25), .B(
        LED_128_Instance_mixcolumns_out[4]), .ZN(
        LED_128_Instance_mixcolumns_out[52]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U39 ( .A(
        LED_128_Instance_mixcolumns_out[23]), .B(
        LED_128_Instance_MCS_Instance_1_n28), .ZN(
        LED_128_Instance_MCS_Instance_1_n25) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U38 ( .A(
        LED_128_Instance_subcells_out[50]), .B(
        LED_128_Instance_mixcolumns_out[39]), .Z(
        LED_128_Instance_MCS_Instance_1_n28) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U37 ( .A(
        LED_128_Instance_MCS_Instance_1_n24), .B(
        LED_128_Instance_MCS_Instance_1_n23), .ZN(
        LED_128_Instance_mixcolumns_out[39]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U36 ( .A(
        LED_128_Instance_subcells_out[51]), .B(
        LED_128_Instance_subcells_out[45]), .ZN(
        LED_128_Instance_MCS_Instance_1_n23) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U35 ( .A(
        LED_128_Instance_mixcolumns_out[22]), .B(
        LED_128_Instance_mixcolumns_out[6]), .Z(
        LED_128_Instance_MCS_Instance_1_n24) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U34 ( .A(
        LED_128_Instance_MCS_Instance_1_n22), .B(
        LED_128_Instance_MCS_Instance_1_n21), .ZN(
        LED_128_Instance_mixcolumns_out[22]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U33 ( .A(
        LED_128_Instance_MCS_Instance_1_n20), .B(
        LED_128_Instance_subcells_out[49]), .ZN(
        LED_128_Instance_MCS_Instance_1_n21) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U32 ( .A(
        LED_128_Instance_mixcolumns_out[5]), .B(
        LED_128_Instance_subcells_out[24]), .Z(
        LED_128_Instance_MCS_Instance_1_n22) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U31 ( .A(
        LED_128_Instance_MCS_Instance_1_n19), .B(
        LED_128_Instance_MCS_Instance_1_n18), .ZN(
        LED_128_Instance_mixcolumns_out[5]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U30 ( .A(
        LED_128_Instance_subcells_out[44]), .B(
        LED_128_Instance_subcells_out[47]), .ZN(
        LED_128_Instance_MCS_Instance_1_n18) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U29 ( .A(
        LED_128_Instance_MCS_Instance_1_n17), .B(
        LED_128_Instance_MCS_Instance_1_n34), .Z(
        LED_128_Instance_MCS_Instance_1_n19) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U28 ( .A(
        LED_128_Instance_MCS_Instance_1_n16), .B(
        LED_128_Instance_subcells_out[6]), .ZN(
        LED_128_Instance_MCS_Instance_1_n34) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U27 ( .A(
        LED_128_Instance_subcells_out[25]), .B(
        LED_128_Instance_subcells_out[7]), .ZN(
        LED_128_Instance_MCS_Instance_1_n16) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U26 ( .A(
        LED_128_Instance_MCS_Instance_1_n15), .B(
        LED_128_Instance_MCS_Instance_1_n31), .ZN(
        LED_128_Instance_mixcolumns_out[37]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U25 ( .A(
        LED_128_Instance_mixcolumns_out[20]), .B(
        LED_128_Instance_mixcolumns_out[23]), .ZN(
        LED_128_Instance_MCS_Instance_1_n31) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U24 ( .A(
        LED_128_Instance_MCS_Instance_1_n14), .B(
        LED_128_Instance_MCS_Instance_1_n13), .ZN(
        LED_128_Instance_MCS_Instance_1_n15) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U23 ( .A(
        LED_128_Instance_subcells_out[46]), .B(
        LED_128_Instance_subcells_out[47]), .ZN(
        LED_128_Instance_MCS_Instance_1_n13) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U22 ( .A(
        LED_128_Instance_MCS_Instance_1_n12), .B(
        LED_128_Instance_subcells_out[49]), .Z(
        LED_128_Instance_MCS_Instance_1_n14) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U21 ( .A(
        LED_128_Instance_MCS_Instance_1_n11), .B(
        LED_128_Instance_MCS_Instance_1_n10), .ZN(
        LED_128_Instance_mixcolumns_out[20]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U20 ( .A(
        LED_128_Instance_mixcolumns_out[7]), .B(
        LED_128_Instance_subcells_out[51]), .ZN(
        LED_128_Instance_MCS_Instance_1_n10) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U19 ( .A(
        LED_128_Instance_subcells_out[44]), .B(
        LED_128_Instance_subcells_out[26]), .Z(
        LED_128_Instance_MCS_Instance_1_n11) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U18 ( .A(
        LED_128_Instance_MCS_Instance_1_n9), .B(
        LED_128_Instance_MCS_Instance_1_n8), .ZN(
        LED_128_Instance_mixcolumns_out[23]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U17 ( .A(
        LED_128_Instance_subcells_out[50]), .B(
        LED_128_Instance_subcells_out[47]), .ZN(
        LED_128_Instance_MCS_Instance_1_n8) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U16 ( .A(
        LED_128_Instance_mixcolumns_out[6]), .B(
        LED_128_Instance_subcells_out[25]), .Z(
        LED_128_Instance_MCS_Instance_1_n9) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U15 ( .A(
        LED_128_Instance_MCS_Instance_1_n7), .B(
        LED_128_Instance_MCS_Instance_1_n6), .ZN(
        LED_128_Instance_mixcolumns_out[6]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U14 ( .A(
        LED_128_Instance_MCS_Instance_1_n5), .B(
        LED_128_Instance_subcells_out[7]), .ZN(
        LED_128_Instance_MCS_Instance_1_n6) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U13 ( .A(
        LED_128_Instance_subcells_out[4]), .B(
        LED_128_Instance_subcells_out[49]), .Z(
        LED_128_Instance_MCS_Instance_1_n7) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U12 ( .A(
        LED_128_Instance_MCS_Instance_1_n17), .B(
        LED_128_Instance_MCS_Instance_1_n35), .Z(
        LED_128_Instance_mixcolumns_out[21]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U11 ( .A(
        LED_128_Instance_MCS_Instance_1_n4), .B(
        LED_128_Instance_MCS_Instance_1_n12), .ZN(
        LED_128_Instance_MCS_Instance_1_n35) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U10 ( .A(
        LED_128_Instance_mixcolumns_out[7]), .B(
        LED_128_Instance_mixcolumns_out[4]), .Z(
        LED_128_Instance_MCS_Instance_1_n12) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U9 ( .A(
        LED_128_Instance_subcells_out[27]), .B(
        LED_128_Instance_MCS_Instance_1_n5), .ZN(
        LED_128_Instance_MCS_Instance_1_n4) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U8 ( .A(
        LED_128_Instance_subcells_out[26]), .B(
        LED_128_Instance_subcells_out[45]), .Z(
        LED_128_Instance_MCS_Instance_1_n5) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U7 ( .A(
        LED_128_Instance_subcells_out[51]), .B(
        LED_128_Instance_subcells_out[48]), .Z(
        LED_128_Instance_MCS_Instance_1_n17) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U6 ( .A(
        LED_128_Instance_MCS_Instance_1_n3), .B(
        LED_128_Instance_MCS_Instance_1_n2), .ZN(
        LED_128_Instance_mixcolumns_out[4]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U5 ( .A(
        LED_128_Instance_subcells_out[51]), .B(
        LED_128_Instance_subcells_out[47]), .ZN(
        LED_128_Instance_MCS_Instance_1_n2) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U4 ( .A(
        LED_128_Instance_subcells_out[6]), .B(
        LED_128_Instance_subcells_out[24]), .Z(
        LED_128_Instance_MCS_Instance_1_n3) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U3 ( .A(
        LED_128_Instance_MCS_Instance_1_n1), .B(
        LED_128_Instance_subcells_out[50]), .ZN(
        LED_128_Instance_mixcolumns_out[7]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_1_U2 ( .A(
        LED_128_Instance_MCS_Instance_1_n20), .B(
        LED_128_Instance_subcells_out[5]), .ZN(
        LED_128_Instance_MCS_Instance_1_n1) );
  XOR2_X1 LED_128_Instance_MCS_Instance_1_U1 ( .A(
        LED_128_Instance_subcells_out[46]), .B(
        LED_128_Instance_subcells_out[27]), .Z(
        LED_128_Instance_MCS_Instance_1_n20) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U54 ( .A(
        LED_128_Instance_MCS_Instance_2_n38), .B(
        LED_128_Instance_MCS_Instance_2_n37), .ZN(
        LED_128_Instance_mixcolumns_out[59]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U53 ( .A(
        LED_128_Instance_mixcolumns_out[11]), .B(
        LED_128_Instance_subcells_out[53]), .ZN(
        LED_128_Instance_MCS_Instance_2_n37) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U52 ( .A(
        LED_128_Instance_mixcolumns_out[42]), .B(
        LED_128_Instance_mixcolumns_out[26]), .Z(
        LED_128_Instance_MCS_Instance_2_n38) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U51 ( .A(
        LED_128_Instance_MCS_Instance_2_n36), .B(
        LED_128_Instance_MCS_Instance_2_n35), .ZN(
        LED_128_Instance_mixcolumns_out[42]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U50 ( .A(
        LED_128_Instance_subcells_out[54]), .B(
        LED_128_Instance_MCS_Instance_2_n34), .ZN(
        LED_128_Instance_MCS_Instance_2_n36) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U49 ( .A(
        LED_128_Instance_MCS_Instance_2_n33), .B(
        LED_128_Instance_mixcolumns_out[41]), .ZN(
        LED_128_Instance_mixcolumns_out[58]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U48 ( .A(
        LED_128_Instance_mixcolumns_out[10]), .B(
        LED_128_Instance_MCS_Instance_2_n35), .ZN(
        LED_128_Instance_MCS_Instance_2_n33) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U47 ( .A(
        LED_128_Instance_MCS_Instance_2_n32), .B(
        LED_128_Instance_MCS_Instance_2_n31), .ZN(
        LED_128_Instance_mixcolumns_out[57]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U46 ( .A(
        LED_128_Instance_MCS_Instance_2_n30), .B(
        LED_128_Instance_MCS_Instance_2_n29), .ZN(
        LED_128_Instance_MCS_Instance_2_n32) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U45 ( .A(
        LED_128_Instance_subcells_out[55]), .B(
        LED_128_Instance_mixcolumns_out[9]), .ZN(
        LED_128_Instance_MCS_Instance_2_n29) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U44 ( .A(
        LED_128_Instance_mixcolumns_out[40]), .B(
        LED_128_Instance_MCS_Instance_2_n28), .Z(
        LED_128_Instance_MCS_Instance_2_n30) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U43 ( .A(
        LED_128_Instance_MCS_Instance_2_n27), .B(
        LED_128_Instance_MCS_Instance_2_n26), .ZN(
        LED_128_Instance_mixcolumns_out[40]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U42 ( .A(
        LED_128_Instance_subcells_out[34]), .B(
        LED_128_Instance_mixcolumns_out[11]), .ZN(
        LED_128_Instance_MCS_Instance_2_n26) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U41 ( .A(
        LED_128_Instance_subcells_out[52]), .B(
        LED_128_Instance_mixcolumns_out[27]), .Z(
        LED_128_Instance_MCS_Instance_2_n27) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U40 ( .A(
        LED_128_Instance_MCS_Instance_2_n25), .B(
        LED_128_Instance_mixcolumns_out[8]), .ZN(
        LED_128_Instance_mixcolumns_out[56]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U39 ( .A(
        LED_128_Instance_mixcolumns_out[27]), .B(
        LED_128_Instance_MCS_Instance_2_n28), .ZN(
        LED_128_Instance_MCS_Instance_2_n25) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U38 ( .A(
        LED_128_Instance_subcells_out[54]), .B(
        LED_128_Instance_mixcolumns_out[43]), .Z(
        LED_128_Instance_MCS_Instance_2_n28) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U37 ( .A(
        LED_128_Instance_MCS_Instance_2_n24), .B(
        LED_128_Instance_MCS_Instance_2_n23), .ZN(
        LED_128_Instance_mixcolumns_out[43]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U36 ( .A(
        LED_128_Instance_subcells_out[55]), .B(
        LED_128_Instance_subcells_out[33]), .ZN(
        LED_128_Instance_MCS_Instance_2_n23) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U35 ( .A(
        LED_128_Instance_mixcolumns_out[26]), .B(
        LED_128_Instance_mixcolumns_out[10]), .Z(
        LED_128_Instance_MCS_Instance_2_n24) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U34 ( .A(
        LED_128_Instance_MCS_Instance_2_n22), .B(
        LED_128_Instance_MCS_Instance_2_n21), .ZN(
        LED_128_Instance_mixcolumns_out[26]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U33 ( .A(
        LED_128_Instance_MCS_Instance_2_n20), .B(
        LED_128_Instance_subcells_out[53]), .ZN(
        LED_128_Instance_MCS_Instance_2_n21) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U32 ( .A(
        LED_128_Instance_mixcolumns_out[9]), .B(
        LED_128_Instance_subcells_out[28]), .Z(
        LED_128_Instance_MCS_Instance_2_n22) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U31 ( .A(
        LED_128_Instance_MCS_Instance_2_n19), .B(
        LED_128_Instance_MCS_Instance_2_n18), .ZN(
        LED_128_Instance_mixcolumns_out[9]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U30 ( .A(
        LED_128_Instance_subcells_out[32]), .B(
        LED_128_Instance_subcells_out[35]), .ZN(
        LED_128_Instance_MCS_Instance_2_n18) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U29 ( .A(
        LED_128_Instance_MCS_Instance_2_n17), .B(
        LED_128_Instance_MCS_Instance_2_n34), .Z(
        LED_128_Instance_MCS_Instance_2_n19) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U28 ( .A(
        LED_128_Instance_MCS_Instance_2_n16), .B(
        LED_128_Instance_subcells_out[10]), .ZN(
        LED_128_Instance_MCS_Instance_2_n34) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U27 ( .A(
        LED_128_Instance_subcells_out[29]), .B(
        LED_128_Instance_subcells_out[11]), .ZN(
        LED_128_Instance_MCS_Instance_2_n16) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U26 ( .A(
        LED_128_Instance_MCS_Instance_2_n15), .B(
        LED_128_Instance_MCS_Instance_2_n31), .ZN(
        LED_128_Instance_mixcolumns_out[41]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U25 ( .A(
        LED_128_Instance_mixcolumns_out[24]), .B(
        LED_128_Instance_mixcolumns_out[27]), .ZN(
        LED_128_Instance_MCS_Instance_2_n31) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U24 ( .A(
        LED_128_Instance_MCS_Instance_2_n14), .B(
        LED_128_Instance_MCS_Instance_2_n13), .ZN(
        LED_128_Instance_MCS_Instance_2_n15) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U23 ( .A(
        LED_128_Instance_subcells_out[34]), .B(
        LED_128_Instance_subcells_out[35]), .ZN(
        LED_128_Instance_MCS_Instance_2_n13) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U22 ( .A(
        LED_128_Instance_MCS_Instance_2_n12), .B(
        LED_128_Instance_subcells_out[53]), .Z(
        LED_128_Instance_MCS_Instance_2_n14) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U21 ( .A(
        LED_128_Instance_MCS_Instance_2_n11), .B(
        LED_128_Instance_MCS_Instance_2_n10), .ZN(
        LED_128_Instance_mixcolumns_out[24]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U20 ( .A(
        LED_128_Instance_mixcolumns_out[11]), .B(
        LED_128_Instance_subcells_out[55]), .ZN(
        LED_128_Instance_MCS_Instance_2_n10) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U19 ( .A(
        LED_128_Instance_subcells_out[32]), .B(
        LED_128_Instance_subcells_out[30]), .Z(
        LED_128_Instance_MCS_Instance_2_n11) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U18 ( .A(
        LED_128_Instance_MCS_Instance_2_n9), .B(
        LED_128_Instance_MCS_Instance_2_n8), .ZN(
        LED_128_Instance_mixcolumns_out[27]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U17 ( .A(
        LED_128_Instance_subcells_out[54]), .B(
        LED_128_Instance_subcells_out[35]), .ZN(
        LED_128_Instance_MCS_Instance_2_n8) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U16 ( .A(
        LED_128_Instance_mixcolumns_out[10]), .B(
        LED_128_Instance_subcells_out[29]), .Z(
        LED_128_Instance_MCS_Instance_2_n9) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U15 ( .A(
        LED_128_Instance_MCS_Instance_2_n7), .B(
        LED_128_Instance_MCS_Instance_2_n6), .ZN(
        LED_128_Instance_mixcolumns_out[10]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U14 ( .A(
        LED_128_Instance_MCS_Instance_2_n5), .B(
        LED_128_Instance_subcells_out[11]), .ZN(
        LED_128_Instance_MCS_Instance_2_n6) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U13 ( .A(
        LED_128_Instance_subcells_out[8]), .B(
        LED_128_Instance_subcells_out[53]), .Z(
        LED_128_Instance_MCS_Instance_2_n7) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U12 ( .A(
        LED_128_Instance_MCS_Instance_2_n17), .B(
        LED_128_Instance_MCS_Instance_2_n35), .Z(
        LED_128_Instance_mixcolumns_out[25]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U11 ( .A(
        LED_128_Instance_MCS_Instance_2_n4), .B(
        LED_128_Instance_MCS_Instance_2_n12), .ZN(
        LED_128_Instance_MCS_Instance_2_n35) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U10 ( .A(
        LED_128_Instance_mixcolumns_out[11]), .B(
        LED_128_Instance_mixcolumns_out[8]), .Z(
        LED_128_Instance_MCS_Instance_2_n12) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U9 ( .A(
        LED_128_Instance_subcells_out[31]), .B(
        LED_128_Instance_MCS_Instance_2_n5), .ZN(
        LED_128_Instance_MCS_Instance_2_n4) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U8 ( .A(
        LED_128_Instance_subcells_out[30]), .B(
        LED_128_Instance_subcells_out[33]), .Z(
        LED_128_Instance_MCS_Instance_2_n5) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U7 ( .A(
        LED_128_Instance_subcells_out[55]), .B(
        LED_128_Instance_subcells_out[52]), .Z(
        LED_128_Instance_MCS_Instance_2_n17) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U6 ( .A(
        LED_128_Instance_MCS_Instance_2_n3), .B(
        LED_128_Instance_MCS_Instance_2_n2), .ZN(
        LED_128_Instance_mixcolumns_out[8]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U5 ( .A(
        LED_128_Instance_subcells_out[55]), .B(
        LED_128_Instance_subcells_out[35]), .ZN(
        LED_128_Instance_MCS_Instance_2_n2) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U4 ( .A(
        LED_128_Instance_subcells_out[10]), .B(
        LED_128_Instance_subcells_out[28]), .Z(
        LED_128_Instance_MCS_Instance_2_n3) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U3 ( .A(
        LED_128_Instance_MCS_Instance_2_n1), .B(
        LED_128_Instance_subcells_out[54]), .ZN(
        LED_128_Instance_mixcolumns_out[11]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_2_U2 ( .A(
        LED_128_Instance_MCS_Instance_2_n20), .B(
        LED_128_Instance_subcells_out[9]), .ZN(
        LED_128_Instance_MCS_Instance_2_n1) );
  XOR2_X1 LED_128_Instance_MCS_Instance_2_U1 ( .A(
        LED_128_Instance_subcells_out[34]), .B(
        LED_128_Instance_subcells_out[31]), .Z(
        LED_128_Instance_MCS_Instance_2_n20) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U54 ( .A(
        LED_128_Instance_MCS_Instance_3_n38), .B(
        LED_128_Instance_MCS_Instance_3_n37), .ZN(
        LED_128_Instance_mixcolumns_out[63]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U53 ( .A(
        LED_128_Instance_mixcolumns_out[15]), .B(
        LED_128_Instance_subcells_out[57]), .ZN(
        LED_128_Instance_MCS_Instance_3_n37) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U52 ( .A(
        LED_128_Instance_mixcolumns_out[46]), .B(
        LED_128_Instance_mixcolumns_out[30]), .Z(
        LED_128_Instance_MCS_Instance_3_n38) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U51 ( .A(
        LED_128_Instance_MCS_Instance_3_n36), .B(
        LED_128_Instance_MCS_Instance_3_n35), .ZN(
        LED_128_Instance_mixcolumns_out[46]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U50 ( .A(
        LED_128_Instance_subcells_out[58]), .B(
        LED_128_Instance_MCS_Instance_3_n34), .ZN(
        LED_128_Instance_MCS_Instance_3_n36) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U49 ( .A(
        LED_128_Instance_MCS_Instance_3_n33), .B(
        LED_128_Instance_mixcolumns_out[45]), .ZN(
        LED_128_Instance_mixcolumns_out[62]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U48 ( .A(
        LED_128_Instance_mixcolumns_out[14]), .B(
        LED_128_Instance_MCS_Instance_3_n35), .ZN(
        LED_128_Instance_MCS_Instance_3_n33) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U47 ( .A(
        LED_128_Instance_MCS_Instance_3_n32), .B(
        LED_128_Instance_MCS_Instance_3_n31), .ZN(
        LED_128_Instance_mixcolumns_out[61]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U46 ( .A(
        LED_128_Instance_MCS_Instance_3_n30), .B(
        LED_128_Instance_MCS_Instance_3_n29), .ZN(
        LED_128_Instance_MCS_Instance_3_n32) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U45 ( .A(
        LED_128_Instance_subcells_out[59]), .B(
        LED_128_Instance_mixcolumns_out[13]), .ZN(
        LED_128_Instance_MCS_Instance_3_n29) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U44 ( .A(
        LED_128_Instance_mixcolumns_out[44]), .B(
        LED_128_Instance_MCS_Instance_3_n28), .Z(
        LED_128_Instance_MCS_Instance_3_n30) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U43 ( .A(
        LED_128_Instance_MCS_Instance_3_n27), .B(
        LED_128_Instance_MCS_Instance_3_n26), .ZN(
        LED_128_Instance_mixcolumns_out[44]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U42 ( .A(
        LED_128_Instance_subcells_out[38]), .B(
        LED_128_Instance_mixcolumns_out[15]), .ZN(
        LED_128_Instance_MCS_Instance_3_n26) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U41 ( .A(
        LED_128_Instance_subcells_out[56]), .B(
        LED_128_Instance_mixcolumns_out[31]), .Z(
        LED_128_Instance_MCS_Instance_3_n27) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U40 ( .A(
        LED_128_Instance_MCS_Instance_3_n25), .B(
        LED_128_Instance_mixcolumns_out[12]), .ZN(
        LED_128_Instance_mixcolumns_out[60]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U39 ( .A(
        LED_128_Instance_mixcolumns_out[31]), .B(
        LED_128_Instance_MCS_Instance_3_n28), .ZN(
        LED_128_Instance_MCS_Instance_3_n25) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U38 ( .A(
        LED_128_Instance_subcells_out[58]), .B(
        LED_128_Instance_mixcolumns_out[47]), .Z(
        LED_128_Instance_MCS_Instance_3_n28) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U37 ( .A(
        LED_128_Instance_MCS_Instance_3_n24), .B(
        LED_128_Instance_MCS_Instance_3_n23), .ZN(
        LED_128_Instance_mixcolumns_out[47]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U36 ( .A(
        LED_128_Instance_subcells_out[59]), .B(
        LED_128_Instance_subcells_out[37]), .ZN(
        LED_128_Instance_MCS_Instance_3_n23) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U35 ( .A(
        LED_128_Instance_mixcolumns_out[30]), .B(
        LED_128_Instance_mixcolumns_out[14]), .Z(
        LED_128_Instance_MCS_Instance_3_n24) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U34 ( .A(
        LED_128_Instance_MCS_Instance_3_n22), .B(
        LED_128_Instance_MCS_Instance_3_n21), .ZN(
        LED_128_Instance_mixcolumns_out[30]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U33 ( .A(
        LED_128_Instance_MCS_Instance_3_n20), .B(
        LED_128_Instance_subcells_out[57]), .ZN(
        LED_128_Instance_MCS_Instance_3_n21) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U32 ( .A(
        LED_128_Instance_mixcolumns_out[13]), .B(
        LED_128_Instance_subcells_out[16]), .Z(
        LED_128_Instance_MCS_Instance_3_n22) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U31 ( .A(
        LED_128_Instance_MCS_Instance_3_n19), .B(
        LED_128_Instance_MCS_Instance_3_n18), .ZN(
        LED_128_Instance_mixcolumns_out[13]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U30 ( .A(
        LED_128_Instance_subcells_out[36]), .B(
        LED_128_Instance_subcells_out[39]), .ZN(
        LED_128_Instance_MCS_Instance_3_n18) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U29 ( .A(
        LED_128_Instance_MCS_Instance_3_n17), .B(
        LED_128_Instance_MCS_Instance_3_n34), .Z(
        LED_128_Instance_MCS_Instance_3_n19) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U28 ( .A(
        LED_128_Instance_MCS_Instance_3_n16), .B(
        LED_128_Instance_subcells_out[14]), .ZN(
        LED_128_Instance_MCS_Instance_3_n34) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U27 ( .A(
        LED_128_Instance_subcells_out[17]), .B(
        LED_128_Instance_subcells_out[15]), .ZN(
        LED_128_Instance_MCS_Instance_3_n16) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U26 ( .A(
        LED_128_Instance_MCS_Instance_3_n15), .B(
        LED_128_Instance_MCS_Instance_3_n31), .ZN(
        LED_128_Instance_mixcolumns_out[45]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U25 ( .A(
        LED_128_Instance_mixcolumns_out[28]), .B(
        LED_128_Instance_mixcolumns_out[31]), .ZN(
        LED_128_Instance_MCS_Instance_3_n31) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U24 ( .A(
        LED_128_Instance_MCS_Instance_3_n14), .B(
        LED_128_Instance_MCS_Instance_3_n13), .ZN(
        LED_128_Instance_MCS_Instance_3_n15) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U23 ( .A(
        LED_128_Instance_subcells_out[38]), .B(
        LED_128_Instance_subcells_out[39]), .ZN(
        LED_128_Instance_MCS_Instance_3_n13) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U22 ( .A(
        LED_128_Instance_MCS_Instance_3_n12), .B(
        LED_128_Instance_subcells_out[57]), .Z(
        LED_128_Instance_MCS_Instance_3_n14) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U21 ( .A(
        LED_128_Instance_MCS_Instance_3_n11), .B(
        LED_128_Instance_MCS_Instance_3_n10), .ZN(
        LED_128_Instance_mixcolumns_out[28]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U20 ( .A(
        LED_128_Instance_mixcolumns_out[15]), .B(
        LED_128_Instance_subcells_out[59]), .ZN(
        LED_128_Instance_MCS_Instance_3_n10) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U19 ( .A(
        LED_128_Instance_subcells_out[36]), .B(
        LED_128_Instance_subcells_out[18]), .Z(
        LED_128_Instance_MCS_Instance_3_n11) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U18 ( .A(
        LED_128_Instance_MCS_Instance_3_n9), .B(
        LED_128_Instance_MCS_Instance_3_n8), .ZN(
        LED_128_Instance_mixcolumns_out[31]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U17 ( .A(
        LED_128_Instance_subcells_out[58]), .B(
        LED_128_Instance_subcells_out[39]), .ZN(
        LED_128_Instance_MCS_Instance_3_n8) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U16 ( .A(
        LED_128_Instance_mixcolumns_out[14]), .B(
        LED_128_Instance_subcells_out[17]), .Z(
        LED_128_Instance_MCS_Instance_3_n9) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U15 ( .A(
        LED_128_Instance_MCS_Instance_3_n7), .B(
        LED_128_Instance_MCS_Instance_3_n6), .ZN(
        LED_128_Instance_mixcolumns_out[14]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U14 ( .A(
        LED_128_Instance_MCS_Instance_3_n5), .B(
        LED_128_Instance_subcells_out[15]), .ZN(
        LED_128_Instance_MCS_Instance_3_n6) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U13 ( .A(
        LED_128_Instance_subcells_out[12]), .B(
        LED_128_Instance_subcells_out[57]), .Z(
        LED_128_Instance_MCS_Instance_3_n7) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U12 ( .A(
        LED_128_Instance_MCS_Instance_3_n17), .B(
        LED_128_Instance_MCS_Instance_3_n35), .Z(
        LED_128_Instance_mixcolumns_out[29]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U11 ( .A(
        LED_128_Instance_MCS_Instance_3_n4), .B(
        LED_128_Instance_MCS_Instance_3_n12), .ZN(
        LED_128_Instance_MCS_Instance_3_n35) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U10 ( .A(
        LED_128_Instance_mixcolumns_out[15]), .B(
        LED_128_Instance_mixcolumns_out[12]), .Z(
        LED_128_Instance_MCS_Instance_3_n12) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U9 ( .A(
        LED_128_Instance_subcells_out[19]), .B(
        LED_128_Instance_MCS_Instance_3_n5), .ZN(
        LED_128_Instance_MCS_Instance_3_n4) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U8 ( .A(
        LED_128_Instance_subcells_out[18]), .B(
        LED_128_Instance_subcells_out[37]), .Z(
        LED_128_Instance_MCS_Instance_3_n5) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U7 ( .A(
        LED_128_Instance_subcells_out[59]), .B(
        LED_128_Instance_subcells_out[56]), .Z(
        LED_128_Instance_MCS_Instance_3_n17) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U6 ( .A(
        LED_128_Instance_MCS_Instance_3_n3), .B(
        LED_128_Instance_MCS_Instance_3_n2), .ZN(
        LED_128_Instance_mixcolumns_out[12]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U5 ( .A(
        LED_128_Instance_subcells_out[59]), .B(
        LED_128_Instance_subcells_out[39]), .ZN(
        LED_128_Instance_MCS_Instance_3_n2) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U4 ( .A(
        LED_128_Instance_subcells_out[14]), .B(
        LED_128_Instance_subcells_out[16]), .Z(
        LED_128_Instance_MCS_Instance_3_n3) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U3 ( .A(
        LED_128_Instance_MCS_Instance_3_n1), .B(
        LED_128_Instance_subcells_out[58]), .ZN(
        LED_128_Instance_mixcolumns_out[15]) );
  XNOR2_X1 LED_128_Instance_MCS_Instance_3_U2 ( .A(
        LED_128_Instance_MCS_Instance_3_n20), .B(
        LED_128_Instance_subcells_out[13]), .ZN(
        LED_128_Instance_MCS_Instance_3_n1) );
  XOR2_X1 LED_128_Instance_MCS_Instance_3_U1 ( .A(
        LED_128_Instance_subcells_out[38]), .B(
        LED_128_Instance_subcells_out[19]), .Z(
        LED_128_Instance_MCS_Instance_3_n20) );
  INV_X1 LED_128_Instance_ks_reg_0__U1 ( .A(LED_128_Instance_ks_reg_0__Q), 
        .ZN(LED_128_Instance_n4) );
  DFF_X1 LED_128_Instance_ks_reg_0__FF_FF ( .D(LED_128_Instance_N10), .CK(CLK), 
        .Q(LED_128_Instance_ks_reg_0__Q), .QN() );
  INV_X1 LED_128_Instance_ks_reg_1__U1 ( .A(LED_128_Instance_n26), .ZN(
        LED_128_Instance_n8) );
  DFF_X1 LED_128_Instance_ks_reg_1__FF_FF ( .D(LED_128_Instance_N11), .CK(CLK), 
        .Q(LED_128_Instance_n26), .QN() );
  INV_X1 LED_128_Instance_ks_reg_2__U1 ( .A(LED_128_Instance_n25), .ZN(
        LED_128_Instance_n1) );
  DFF_X1 LED_128_Instance_ks_reg_2__FF_FF ( .D(LED_128_Instance_N12), .CK(CLK), 
        .Q(LED_128_Instance_n25), .QN() );
  INV_X1 LED_128_Instance_ks_reg_3__U1 ( .A(LED_128_Instance_n2), .ZN(
        LED_128_Instance_n24) );
  DFF_X1 LED_128_Instance_ks_reg_3__FF_FF ( .D(LED_128_Instance_N13), .CK(CLK), 
        .Q(LED_128_Instance_n2), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_0__U1 ( .A(roundconstant[0]), .ZN(
        LED_128_Instance_n6) );
  DFF_X1 LED_128_Instance_roundconstant_reg_0__FF_FF ( .D(LED_128_Instance_N4), 
        .CK(CLK), .Q(roundconstant[0]), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_1__U1 ( .A(roundconstant[1]), .ZN(
        LED_128_Instance_n29) );
  DFF_X1 LED_128_Instance_roundconstant_reg_1__FF_FF ( .D(LED_128_Instance_N5), 
        .CK(CLK), .Q(roundconstant[1]), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_2__U1 ( .A(roundconstant[2]), .ZN(
        LED_128_Instance_n5) );
  DFF_X1 LED_128_Instance_roundconstant_reg_2__FF_FF ( .D(LED_128_Instance_N6), 
        .CK(CLK), .Q(roundconstant[2]), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_3__U1 ( .A(roundconstant[3]), .ZN(
        LED_128_Instance_n30) );
  DFF_X1 LED_128_Instance_roundconstant_reg_3__FF_FF ( .D(LED_128_Instance_N7), 
        .CK(CLK), .Q(roundconstant[3]), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_4__U1 ( .A(roundconstant[4]), .ZN(
        LED_128_Instance_n28) );
  DFF_X1 LED_128_Instance_roundconstant_reg_4__FF_FF ( .D(LED_128_Instance_N8), 
        .CK(CLK), .Q(roundconstant[4]), .QN() );
  INV_X1 LED_128_Instance_roundconstant_reg_5__U1 ( .A(roundconstant[5]), .ZN(
        LED_128_Instance_n27) );
  DFF_X1 LED_128_Instance_roundconstant_reg_5__FF_FF ( .D(LED_128_Instance_N9), 
        .CK(CLK), .Q(roundconstant[5]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_0__U1 ( .A(OUT_ciphertext[0]), .ZN(
        LED_128_Instance_cipherstate_reg_0__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_0__FF_FF ( .D(
        LED_128_Instance_state1[0]), .CK(CLK), .Q(OUT_ciphertext[0]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_1__U1 ( .A(OUT_ciphertext[1]), .ZN(
        LED_128_Instance_cipherstate_reg_1__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_1__FF_FF ( .D(
        LED_128_Instance_state1[1]), .CK(CLK), .Q(OUT_ciphertext[1]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_2__U1 ( .A(OUT_ciphertext[2]), .ZN(
        LED_128_Instance_cipherstate_reg_2__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_2__FF_FF ( .D(
        LED_128_Instance_state1[2]), .CK(CLK), .Q(OUT_ciphertext[2]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_3__U1 ( .A(OUT_ciphertext[3]), .ZN(
        LED_128_Instance_cipherstate_reg_3__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_3__FF_FF ( .D(
        LED_128_Instance_state1[3]), .CK(CLK), .Q(OUT_ciphertext[3]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_4__U1 ( .A(OUT_ciphertext[4]), .ZN(
        LED_128_Instance_cipherstate_reg_4__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_4__FF_FF ( .D(
        LED_128_Instance_state1[4]), .CK(CLK), .Q(OUT_ciphertext[4]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_5__U1 ( .A(OUT_ciphertext[5]), .ZN(
        LED_128_Instance_cipherstate_reg_5__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_5__FF_FF ( .D(
        LED_128_Instance_state1[5]), .CK(CLK), .Q(OUT_ciphertext[5]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_6__U1 ( .A(OUT_ciphertext[6]), .ZN(
        LED_128_Instance_cipherstate_reg_6__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_6__FF_FF ( .D(
        LED_128_Instance_state1[6]), .CK(CLK), .Q(OUT_ciphertext[6]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_7__U1 ( .A(OUT_ciphertext[7]), .ZN(
        LED_128_Instance_cipherstate_reg_7__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_7__FF_FF ( .D(
        LED_128_Instance_state1[7]), .CK(CLK), .Q(OUT_ciphertext[7]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_8__U1 ( .A(OUT_ciphertext[8]), .ZN(
        LED_128_Instance_cipherstate_reg_8__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_8__FF_FF ( .D(
        LED_128_Instance_state1[8]), .CK(CLK), .Q(OUT_ciphertext[8]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_9__U1 ( .A(OUT_ciphertext[9]), .ZN(
        LED_128_Instance_cipherstate_reg_9__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_9__FF_FF ( .D(
        LED_128_Instance_state1[9]), .CK(CLK), .Q(OUT_ciphertext[9]), .QN() );
  INV_X1 LED_128_Instance_cipherstate_reg_10__U1 ( .A(OUT_ciphertext[10]), 
        .ZN(LED_128_Instance_cipherstate_reg_10__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_10__FF_FF ( .D(
        LED_128_Instance_state1[10]), .CK(CLK), .Q(OUT_ciphertext[10]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_11__U1 ( .A(OUT_ciphertext[11]), 
        .ZN(LED_128_Instance_cipherstate_reg_11__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_11__FF_FF ( .D(
        LED_128_Instance_state1[11]), .CK(CLK), .Q(OUT_ciphertext[11]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_12__U1 ( .A(OUT_ciphertext[12]), 
        .ZN(LED_128_Instance_cipherstate_reg_12__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_12__FF_FF ( .D(
        LED_128_Instance_state1[12]), .CK(CLK), .Q(OUT_ciphertext[12]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_13__U1 ( .A(OUT_ciphertext[13]), 
        .ZN(LED_128_Instance_cipherstate_reg_13__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_13__FF_FF ( .D(
        LED_128_Instance_state1[13]), .CK(CLK), .Q(OUT_ciphertext[13]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_14__U1 ( .A(OUT_ciphertext[14]), 
        .ZN(LED_128_Instance_cipherstate_reg_14__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_14__FF_FF ( .D(
        LED_128_Instance_state1[14]), .CK(CLK), .Q(OUT_ciphertext[14]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_15__U1 ( .A(OUT_ciphertext[15]), 
        .ZN(LED_128_Instance_cipherstate_reg_15__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_15__FF_FF ( .D(
        LED_128_Instance_state1[15]), .CK(CLK), .Q(OUT_ciphertext[15]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_16__U1 ( .A(OUT_ciphertext[16]), 
        .ZN(LED_128_Instance_cipherstate_reg_16__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_16__FF_FF ( .D(
        LED_128_Instance_state1[16]), .CK(CLK), .Q(OUT_ciphertext[16]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_17__U1 ( .A(OUT_ciphertext[17]), 
        .ZN(LED_128_Instance_cipherstate_reg_17__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_17__FF_FF ( .D(
        LED_128_Instance_state1[17]), .CK(CLK), .Q(OUT_ciphertext[17]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_18__U1 ( .A(OUT_ciphertext[18]), 
        .ZN(LED_128_Instance_cipherstate_reg_18__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_18__FF_FF ( .D(
        LED_128_Instance_state1[18]), .CK(CLK), .Q(OUT_ciphertext[18]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_19__U1 ( .A(OUT_ciphertext[19]), 
        .ZN(LED_128_Instance_cipherstate_reg_19__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_19__FF_FF ( .D(
        LED_128_Instance_state1[19]), .CK(CLK), .Q(OUT_ciphertext[19]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_20__U1 ( .A(OUT_ciphertext[20]), 
        .ZN(LED_128_Instance_cipherstate_reg_20__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_20__FF_FF ( .D(
        LED_128_Instance_state1[20]), .CK(CLK), .Q(OUT_ciphertext[20]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_21__U1 ( .A(OUT_ciphertext[21]), 
        .ZN(LED_128_Instance_cipherstate_reg_21__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_21__FF_FF ( .D(
        LED_128_Instance_state1[21]), .CK(CLK), .Q(OUT_ciphertext[21]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_22__U1 ( .A(OUT_ciphertext[22]), 
        .ZN(LED_128_Instance_cipherstate_reg_22__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_22__FF_FF ( .D(
        LED_128_Instance_state1[22]), .CK(CLK), .Q(OUT_ciphertext[22]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_23__U1 ( .A(OUT_ciphertext[23]), 
        .ZN(LED_128_Instance_cipherstate_reg_23__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_23__FF_FF ( .D(
        LED_128_Instance_state1[23]), .CK(CLK), .Q(OUT_ciphertext[23]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_24__U1 ( .A(OUT_ciphertext[24]), 
        .ZN(LED_128_Instance_cipherstate_reg_24__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_24__FF_FF ( .D(
        LED_128_Instance_state1[24]), .CK(CLK), .Q(OUT_ciphertext[24]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_25__U1 ( .A(OUT_ciphertext[25]), 
        .ZN(LED_128_Instance_cipherstate_reg_25__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_25__FF_FF ( .D(
        LED_128_Instance_state1[25]), .CK(CLK), .Q(OUT_ciphertext[25]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_26__U1 ( .A(OUT_ciphertext[26]), 
        .ZN(LED_128_Instance_cipherstate_reg_26__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_26__FF_FF ( .D(
        LED_128_Instance_state1[26]), .CK(CLK), .Q(OUT_ciphertext[26]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_27__U1 ( .A(OUT_ciphertext[27]), 
        .ZN(LED_128_Instance_cipherstate_reg_27__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_27__FF_FF ( .D(
        LED_128_Instance_state1[27]), .CK(CLK), .Q(OUT_ciphertext[27]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_28__U1 ( .A(OUT_ciphertext[28]), 
        .ZN(LED_128_Instance_cipherstate_reg_28__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_28__FF_FF ( .D(
        LED_128_Instance_state1[28]), .CK(CLK), .Q(OUT_ciphertext[28]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_29__U1 ( .A(OUT_ciphertext[29]), 
        .ZN(LED_128_Instance_cipherstate_reg_29__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_29__FF_FF ( .D(
        LED_128_Instance_state1[29]), .CK(CLK), .Q(OUT_ciphertext[29]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_30__U1 ( .A(OUT_ciphertext[30]), 
        .ZN(LED_128_Instance_cipherstate_reg_30__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_30__FF_FF ( .D(
        LED_128_Instance_state1[30]), .CK(CLK), .Q(OUT_ciphertext[30]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_31__U1 ( .A(OUT_ciphertext[31]), 
        .ZN(LED_128_Instance_cipherstate_reg_31__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_31__FF_FF ( .D(
        LED_128_Instance_state1[31]), .CK(CLK), .Q(OUT_ciphertext[31]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_32__U1 ( .A(OUT_ciphertext[32]), 
        .ZN(LED_128_Instance_cipherstate_reg_32__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_32__FF_FF ( .D(
        LED_128_Instance_state1[32]), .CK(CLK), .Q(OUT_ciphertext[32]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_33__U1 ( .A(OUT_ciphertext[33]), 
        .ZN(LED_128_Instance_cipherstate_reg_33__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_33__FF_FF ( .D(
        LED_128_Instance_state1[33]), .CK(CLK), .Q(OUT_ciphertext[33]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_34__U1 ( .A(OUT_ciphertext[34]), 
        .ZN(LED_128_Instance_cipherstate_reg_34__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_34__FF_FF ( .D(
        LED_128_Instance_state1[34]), .CK(CLK), .Q(OUT_ciphertext[34]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_35__U1 ( .A(OUT_ciphertext[35]), 
        .ZN(LED_128_Instance_cipherstate_reg_35__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_35__FF_FF ( .D(
        LED_128_Instance_state1[35]), .CK(CLK), .Q(OUT_ciphertext[35]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_36__U1 ( .A(OUT_ciphertext[36]), 
        .ZN(LED_128_Instance_cipherstate_reg_36__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_36__FF_FF ( .D(
        LED_128_Instance_state1[36]), .CK(CLK), .Q(OUT_ciphertext[36]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_37__U1 ( .A(OUT_ciphertext[37]), 
        .ZN(LED_128_Instance_cipherstate_reg_37__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_37__FF_FF ( .D(
        LED_128_Instance_state1[37]), .CK(CLK), .Q(OUT_ciphertext[37]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_38__U1 ( .A(OUT_ciphertext[38]), 
        .ZN(LED_128_Instance_cipherstate_reg_38__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_38__FF_FF ( .D(
        LED_128_Instance_state1[38]), .CK(CLK), .Q(OUT_ciphertext[38]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_39__U1 ( .A(OUT_ciphertext[39]), 
        .ZN(LED_128_Instance_cipherstate_reg_39__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_39__FF_FF ( .D(
        LED_128_Instance_state1[39]), .CK(CLK), .Q(OUT_ciphertext[39]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_40__U1 ( .A(OUT_ciphertext[40]), 
        .ZN(LED_128_Instance_cipherstate_reg_40__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_40__FF_FF ( .D(
        LED_128_Instance_state1[40]), .CK(CLK), .Q(OUT_ciphertext[40]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_41__U1 ( .A(OUT_ciphertext[41]), 
        .ZN(LED_128_Instance_cipherstate_reg_41__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_41__FF_FF ( .D(
        LED_128_Instance_state1[41]), .CK(CLK), .Q(OUT_ciphertext[41]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_42__U1 ( .A(OUT_ciphertext[42]), 
        .ZN(LED_128_Instance_cipherstate_reg_42__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_42__FF_FF ( .D(
        LED_128_Instance_state1[42]), .CK(CLK), .Q(OUT_ciphertext[42]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_43__U1 ( .A(OUT_ciphertext[43]), 
        .ZN(LED_128_Instance_cipherstate_reg_43__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_43__FF_FF ( .D(
        LED_128_Instance_state1[43]), .CK(CLK), .Q(OUT_ciphertext[43]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_44__U1 ( .A(OUT_ciphertext[44]), 
        .ZN(LED_128_Instance_cipherstate_reg_44__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_44__FF_FF ( .D(
        LED_128_Instance_state1[44]), .CK(CLK), .Q(OUT_ciphertext[44]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_45__U1 ( .A(OUT_ciphertext[45]), 
        .ZN(LED_128_Instance_cipherstate_reg_45__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_45__FF_FF ( .D(
        LED_128_Instance_state1[45]), .CK(CLK), .Q(OUT_ciphertext[45]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_46__U1 ( .A(OUT_ciphertext[46]), 
        .ZN(LED_128_Instance_cipherstate_reg_46__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_46__FF_FF ( .D(
        LED_128_Instance_state1[46]), .CK(CLK), .Q(OUT_ciphertext[46]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_47__U1 ( .A(OUT_ciphertext[47]), 
        .ZN(LED_128_Instance_cipherstate_reg_47__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_47__FF_FF ( .D(
        LED_128_Instance_state1[47]), .CK(CLK), .Q(OUT_ciphertext[47]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_48__U1 ( .A(OUT_ciphertext[48]), 
        .ZN(LED_128_Instance_cipherstate_reg_48__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_48__FF_FF ( .D(
        LED_128_Instance_state1[48]), .CK(CLK), .Q(OUT_ciphertext[48]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_49__U1 ( .A(OUT_ciphertext[49]), 
        .ZN(LED_128_Instance_cipherstate_reg_49__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_49__FF_FF ( .D(
        LED_128_Instance_state1[49]), .CK(CLK), .Q(OUT_ciphertext[49]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_50__U1 ( .A(OUT_ciphertext[50]), 
        .ZN(LED_128_Instance_cipherstate_reg_50__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_50__FF_FF ( .D(
        LED_128_Instance_state1[50]), .CK(CLK), .Q(OUT_ciphertext[50]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_51__U1 ( .A(OUT_ciphertext[51]), 
        .ZN(LED_128_Instance_cipherstate_reg_51__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_51__FF_FF ( .D(
        LED_128_Instance_state1[51]), .CK(CLK), .Q(OUT_ciphertext[51]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_52__U1 ( .A(OUT_ciphertext[52]), 
        .ZN(LED_128_Instance_cipherstate_reg_52__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_52__FF_FF ( .D(
        LED_128_Instance_state1[52]), .CK(CLK), .Q(OUT_ciphertext[52]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_53__U1 ( .A(OUT_ciphertext[53]), 
        .ZN(LED_128_Instance_cipherstate_reg_53__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_53__FF_FF ( .D(
        LED_128_Instance_state1[53]), .CK(CLK), .Q(OUT_ciphertext[53]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_54__U1 ( .A(OUT_ciphertext[54]), 
        .ZN(LED_128_Instance_cipherstate_reg_54__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_54__FF_FF ( .D(
        LED_128_Instance_state1[54]), .CK(CLK), .Q(OUT_ciphertext[54]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_55__U1 ( .A(OUT_ciphertext[55]), 
        .ZN(LED_128_Instance_cipherstate_reg_55__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_55__FF_FF ( .D(
        LED_128_Instance_state1[55]), .CK(CLK), .Q(OUT_ciphertext[55]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_56__U1 ( .A(OUT_ciphertext[56]), 
        .ZN(LED_128_Instance_cipherstate_reg_56__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_56__FF_FF ( .D(
        LED_128_Instance_state1[56]), .CK(CLK), .Q(OUT_ciphertext[56]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_57__U1 ( .A(OUT_ciphertext[57]), 
        .ZN(LED_128_Instance_cipherstate_reg_57__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_57__FF_FF ( .D(
        LED_128_Instance_state1[57]), .CK(CLK), .Q(OUT_ciphertext[57]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_58__U1 ( .A(OUT_ciphertext[58]), 
        .ZN(LED_128_Instance_cipherstate_reg_58__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_58__FF_FF ( .D(
        LED_128_Instance_state1[58]), .CK(CLK), .Q(OUT_ciphertext[58]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_59__U1 ( .A(OUT_ciphertext[59]), 
        .ZN(LED_128_Instance_cipherstate_reg_59__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_59__FF_FF ( .D(
        LED_128_Instance_state1[59]), .CK(CLK), .Q(OUT_ciphertext[59]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_60__U1 ( .A(OUT_ciphertext[60]), 
        .ZN(LED_128_Instance_cipherstate_reg_60__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_60__FF_FF ( .D(
        LED_128_Instance_state1[60]), .CK(CLK), .Q(OUT_ciphertext[60]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_61__U1 ( .A(OUT_ciphertext[61]), 
        .ZN(LED_128_Instance_cipherstate_reg_61__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_61__FF_FF ( .D(
        LED_128_Instance_state1[61]), .CK(CLK), .Q(OUT_ciphertext[61]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_62__U1 ( .A(OUT_ciphertext[62]), 
        .ZN(LED_128_Instance_cipherstate_reg_62__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_62__FF_FF ( .D(
        LED_128_Instance_state1[62]), .CK(CLK), .Q(OUT_ciphertext[62]), .QN()
         );
  INV_X1 LED_128_Instance_cipherstate_reg_63__U1 ( .A(OUT_ciphertext[63]), 
        .ZN(LED_128_Instance_cipherstate_reg_63__QN) );
  DFF_X1 LED_128_Instance_cipherstate_reg_63__FF_FF ( .D(
        LED_128_Instance_state1[63]), .CK(CLK), .Q(OUT_ciphertext[63]), .QN()
         );
  INV_X1 internal_done_reg_U1 ( .A(OUT_done), .ZN(internal_done_reg_QN) );
  DFF_X1 internal_done_reg_FF_FF ( .D(n15), .CK(CLK), .Q(OUT_done), .QN() );
endmodule

